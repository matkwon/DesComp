library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 16;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant ANDD : std_logic_vector(3 downto 0) := "0100";
  constant LDI  : std_logic_vector(3 downto 0) := "0101";
  constant STA  : std_logic_vector(3 downto 0) := "0110";
  constant JMP  : std_logic_vector(3 downto 0) := "0111";
  constant JEQ  : std_logic_vector(3 downto 0) := "1000";
  constant CEQ  : std_logic_vector(3 downto 0) := "1001";
  constant JSR  : std_logic_vector(3 downto 0) := "1010";
  constant RET  : std_logic_vector(3 downto 0) := "1011";
  constant JNE  : std_logic_vector(3 downto 0) := "1100";
  constant JLT  : std_logic_vector(3 downto 0) := "1101";
  constant CLT  : std_logic_vector(3 downto 0) := "1110";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
  

-- LABEL Setup
tmp(0) := "0101" & "000" & "010000000" ;	-- LDI R0, $128
tmp(1) := "0110" & "000" & "000111111" ;	-- STA @63, R0
tmp(2) := "0101" & "000" & "000000000" ;	-- LDI R0, $0
tmp(3) := "0110" & "000" & "000000000" ;	-- STA @0, R0
tmp(4) := "0101" & "001" & "000000001" ;	-- LDI R1, $1
tmp(5) := "0110" & "001" & "000000001" ;	-- STA @1, R1
tmp(6) := "0101" & "001" & "000000010" ;	-- LDI R1, $2
tmp(7) := "0110" & "001" & "000000010" ;	-- STA @2, R1
tmp(8) := "0101" & "001" & "000000011" ;	-- LDI R1, $3
tmp(9) := "0110" & "001" & "000000011" ;	-- STA @3, R1
tmp(10) := "0110" & "001" & "000010011" ;	-- STA @BAS5, R1
tmp(11) := "0101" & "001" & "000000100" ;	-- LDI R1, $4
tmp(12) := "0110" & "001" & "000000100" ;	-- STA @4, R1
tmp(13) := "0101" & "001" & "000000101" ;	-- LDI R1, $5
tmp(14) := "0110" & "001" & "000000101" ;	-- STA @5, R1
tmp(15) := "0101" & "001" & "000000110" ;	-- LDI R1, $6
tmp(16) := "0110" & "001" & "000000110" ;	-- STA @6, R1
tmp(17) := "0101" & "001" & "000001000" ;	-- LDI R1, $8
tmp(18) := "0110" & "001" & "000001000" ;	-- STA @8, R1
tmp(19) := "0101" & "001" & "000001010" ;	-- LDI R1, $10
tmp(20) := "0110" & "001" & "000001010" ;	-- STA @10, R1
tmp(21) := "0110" & "001" & "000010010" ;	-- STA @BAS4, R1
tmp(22) := "0110" & "000" & "000010001" ;	-- STA @AMPM, R0
tmp(23) := "0110" & "000" & "000001011" ;	-- STA @MEM0, R0
tmp(24) := "0110" & "000" & "000001101" ;	-- STA @MEM2, R0
tmp(25) := "0110" & "000" & "000001100" ;	-- STA @MEM1, R0
tmp(26) := "0110" & "000" & "000001110" ;	-- STA @MEM3, R0
tmp(27) := "0110" & "000" & "000001111" ;	-- STA @MEM4, R0
tmp(28) := "0110" & "000" & "000010000" ;	-- STA @MEM5, R0
tmp(29) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(30) := "0110" & "000" & "100100001" ;	-- STA @HEX1, R0
tmp(31) := "0110" & "000" & "100100010" ;	-- STA @HEX2, R0
tmp(32) := "0110" & "000" & "100100011" ;	-- STA @HEX3, R0
tmp(33) := "0110" & "000" & "100100100" ;	-- STA @HEX4, R0
tmp(34) := "0110" & "000" & "100100101" ;	-- STA @HEX5, R0
tmp(35) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(36) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(37) := "0001" & "101" & "000000000" ;	-- LDA R5, @0
tmp(38) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(39) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(40) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(41) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(42) := "0001" & "000" & "000000000" ;	-- LDA R0, @0

-- LABEL Clock
tmp(43) := "0001" & "011" & "000001011" ;	-- LDA R3, @MEM0
tmp(44) := "0110" & "011" & "100100000" ;	-- STA @HEX0, R3
tmp(45) := "0001" & "011" & "000001100" ;	-- LDA R3, @MEM1
tmp(46) := "0110" & "011" & "100100001" ;	-- STA @HEX1, R3
tmp(47) := "0001" & "011" & "000001101" ;	-- LDA R3, @MEM2
tmp(48) := "0110" & "011" & "100100010" ;	-- STA @HEX2, R3
tmp(49) := "0001" & "011" & "000001110" ;	-- LDA R3, @MEM3
tmp(50) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(51) := "0001" & "011" & "000001111" ;	-- LDA R3, @MEM4
tmp(52) := "0110" & "011" & "100100100" ;	-- STA @HEX4, R3
tmp(53) := "0001" & "011" & "000010000" ;	-- LDA R3, @MEM5
tmp(54) := "0110" & "011" & "100100101" ;	-- STA @HEX5, R3
tmp(55) := "0111" & "000" & "010101101" ;	-- JMP @WaitSet

-- LABEL IncClk
tmp(56) := "0001" & "111" & "101100101" ;	-- LDA R7, @SEC
tmp(57) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(58) := "1001" & "111" & "000000001" ;	-- CEQ R7, @1
tmp(59) := "1100" & "000" & "010101101" ;	-- JNE @WaitSet
tmp(60) := "0110" & "000" & "111111010" ;	-- CLR @SEC
tmp(61) := "0001" & "000" & "000001011" ;	-- LDA R0, @MEM0
tmp(62) := "0010" & "000" & "000000001" ;	-- SOMA R0, @1
tmp(63) := "1001" & "000" & "000001010" ;	-- CEQ R0, @10
tmp(64) := "1000" & "000" & "001000011" ;	-- JEQ @ResetMem0
tmp(65) := "0110" & "000" & "000001011" ;	-- STA @MEM0, R0
tmp(66) := "0111" & "000" & "010101101" ;	-- JMP @WaitSet

-- LABEL ResetMem0
tmp(67) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(68) := "0110" & "000" & "000001011" ;	-- STA @MEM0, R0
tmp(69) := "0001" & "001" & "000001100" ;	-- LDA R1, @MEM1
tmp(70) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(71) := "1001" & "001" & "000000110" ;	-- CEQ R1, @6
tmp(72) := "1000" & "000" & "001001011" ;	-- JEQ @ResetMem1
tmp(73) := "0110" & "001" & "000001100" ;	-- STA @MEM1, R1
tmp(74) := "0111" & "000" & "010101101" ;	-- JMP @WaitSet

-- LABEL ResetMem1
tmp(75) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(76) := "0110" & "001" & "000001100" ;	-- STA @MEM1, R1
tmp(77) := "0001" & "010" & "000001101" ;	-- LDA R2, @MEM2
tmp(78) := "0010" & "010" & "000000001" ;	-- SOMA R2, @1
tmp(79) := "1001" & "010" & "000001010" ;	-- CEQ R2, @10
tmp(80) := "1000" & "000" & "001010011" ;	-- JEQ @ResetMem2
tmp(81) := "0110" & "010" & "000001101" ;	-- STA @MEM2, R2
tmp(82) := "0111" & "000" & "010101101" ;	-- JMP @WaitSet

-- LABEL ResetMem2
tmp(83) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(84) := "0110" & "010" & "000001101" ;	-- STA @MEM2, R2
tmp(85) := "0001" & "011" & "000001110" ;	-- LDA R3, @MEM3
tmp(86) := "0010" & "011" & "000000001" ;	-- SOMA R3, @1
tmp(87) := "1001" & "011" & "000000110" ;	-- CEQ R3, @6
tmp(88) := "1000" & "000" & "001011011" ;	-- JEQ @ResetMem3
tmp(89) := "0110" & "011" & "000001110" ;	-- STA @MEM3, R3
tmp(90) := "0111" & "000" & "010101101" ;	-- JMP @WaitSet

-- LABEL ResetMem3
tmp(91) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(92) := "0110" & "011" & "000001110" ;	-- STA @MEM3, R3
tmp(93) := "0001" & "100" & "000001111" ;	-- LDA R4, @MEM4
tmp(94) := "0010" & "100" & "000000001" ;	-- SOMA R4, @1
tmp(95) := "1001" & "100" & "000010010" ;	-- CEQ R4, @BAS4
tmp(96) := "1000" & "000" & "001100011" ;	-- JEQ @ResetMem4
tmp(97) := "0110" & "100" & "000001111" ;	-- STA @MEM4, R4
tmp(98) := "0111" & "000" & "010101101" ;	-- JMP @WaitSet

-- LABEL ResetMem4
tmp(99) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(100) := "0110" & "100" & "000001111" ;	-- STA @MEM4, R4
tmp(101) := "0001" & "101" & "000010000" ;	-- LDA R5, @MEM5
tmp(102) := "0010" & "101" & "000000001" ;	-- SOMA R5, @1
tmp(103) := "1001" & "101" & "000010011" ;	-- CEQ R5, @BAS5
tmp(104) := "1000" & "000" & "010011110" ;	-- JEQ @Zera
tmp(105) := "0110" & "101" & "000010000" ;	-- STA @MEM5, R5
tmp(106) := "1001" & "101" & "000000010" ;	-- CEQ R5, @2
tmp(107) := "1100" & "000" & "010101101" ;	-- JNE @WaitSet
tmp(108) := "1010" & "000" & "010010010" ;	-- JSR @BAS4SET4
tmp(109) := "0111" & "000" & "010101101" ;	-- JMP @WaitSet

-- LABEL Base12
tmp(110) := "0001" & "101" & "000010000" ;	-- LDA R5, @MEM5
tmp(111) := "0001" & "100" & "000001111" ;	-- LDA R4, @MEM4
tmp(112) := "1001" & "101" & "000000000" ;	-- CEQ R5, @0
tmp(113) := "1000" & "000" & "001111010" ;	-- JEQ @Display4Base12
tmp(114) := "1001" & "101" & "000000001" ;	-- CEQ R5, @1
tmp(115) := "1000" & "000" & "001110111" ;	-- JEQ @VerificaMem4
tmp(116) := "1110" & "100" & "000000010" ;	-- CLT R4, @2
tmp(117) := "1101" & "000" & "010000100" ;	-- JLT @Caso2
tmp(118) := "0111" & "000" & "001111110" ;	-- JMP @Caso1

-- LABEL VerificaMem4
tmp(119) := "1110" & "100" & "000000010" ;	-- CLT R4, @2
tmp(120) := "1101" & "000" & "001111010" ;	-- JLT @Display4Base12
tmp(121) := "0111" & "000" & "001111110" ;	-- JMP @Caso1

-- LABEL Display4Base12
tmp(122) := "0110" & "100" & "100100100" ;	-- STA @HEX4, R4
tmp(123) := "0110" & "101" & "100100101" ;	-- STA @HEX5, R5
tmp(124) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(125) := "0111" & "000" & "010001001" ;	-- JMP @RetConv

-- LABEL Caso1
tmp(126) := "0011" & "100" & "000000010" ;	-- SUB R4, @2
tmp(127) := "0110" & "100" & "100100100" ;	-- STA @HEX4, R4
tmp(128) := "0011" & "101" & "000000001" ;	-- SUB R5, @1
tmp(129) := "0110" & "101" & "100100101" ;	-- STA @HEX5, R5
tmp(130) := "0001" & "111" & "000000001" ;	-- LDA R7, @1
tmp(131) := "0111" & "000" & "010001001" ;	-- JMP @RetConv

-- LABEL Caso2
tmp(132) := "0010" & "100" & "000001000" ;	-- SOMA R4, @8
tmp(133) := "0110" & "100" & "100100100" ;	-- STA @HEX4, R4
tmp(134) := "0011" & "101" & "000000010" ;	-- SUB R5, @2
tmp(135) := "0110" & "101" & "100100101" ;	-- STA @HEX5, R5
tmp(136) := "0001" & "111" & "000000001" ;	-- LDA R7, @1

-- LABEL RetConv
tmp(137) := "0110" & "111" & "100000010" ;	-- STA @LED9, R7
tmp(138) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Base24
tmp(139) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(140) := "0110" & "111" & "100000010" ;	-- STA @LED9, R7
tmp(141) := "0001" & "100" & "000001111" ;	-- LDA R4, @MEM4
tmp(142) := "0110" & "100" & "100100100" ;	-- STA @HEX4, R4
tmp(143) := "0001" & "101" & "000010000" ;	-- LDA R5, @MEM5
tmp(144) := "0110" & "101" & "100100101" ;	-- STA @HEX5, R5
tmp(145) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL BAS4SET4
tmp(146) := "0001" & "100" & "000000100" ;	-- LDA R4, @4
tmp(147) := "0110" & "100" & "000010010" ;	-- STA @BAS4, R4
tmp(148) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL BAS4SET10
tmp(149) := "0001" & "100" & "000001010" ;	-- LDA R4, @10
tmp(150) := "0110" & "100" & "000010010" ;	-- STA @BAS4, R4
tmp(151) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL BAS5SET2
tmp(152) := "0001" & "100" & "000000010" ;	-- LDA R4, @2
tmp(153) := "0110" & "100" & "000010011" ;	-- STA @BAS5, R4
tmp(154) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL BAS5SET3
tmp(155) := "0001" & "100" & "000000011" ;	-- LDA R4, @3
tmp(156) := "0110" & "100" & "000010011" ;	-- STA @BAS5, R4
tmp(157) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Zera
tmp(158) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(159) := "0110" & "000" & "000001011" ;	-- STA @MEM0, R0
tmp(160) := "0110" & "000" & "000001101" ;	-- STA @MEM2, R0
tmp(161) := "0110" & "000" & "000001100" ;	-- STA @MEM1, R0
tmp(162) := "0110" & "000" & "000001110" ;	-- STA @MEM3, R0
tmp(163) := "0110" & "000" & "000001111" ;	-- STA @MEM4, R0
tmp(164) := "0110" & "000" & "000010000" ;	-- STA @MEM5, R0
tmp(165) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(166) := "0110" & "000" & "100100001" ;	-- STA @HEX1, R0
tmp(167) := "0110" & "000" & "100100010" ;	-- STA @HEX2, R0
tmp(168) := "0110" & "000" & "100100011" ;	-- STA @HEX3, R0
tmp(169) := "0110" & "000" & "100100100" ;	-- STA @HEX4, R0
tmp(170) := "0110" & "000" & "100100101" ;	-- STA @HEX5, R0
tmp(171) := "1010" & "000" & "010010101" ;	-- JSR @BAS4SET10
tmp(172) := "0111" & "000" & "010101101" ;	-- JMP @WaitSet

-- LABEL WaitSet
tmp(173) := "0001" & "111" & "101100011" ;	-- LDA R7, @KEY3
tmp(174) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(175) := "1001" & "111" & "000000001" ;	-- CEQ R7, @1
tmp(176) := "1000" & "000" & "011001100" ;	-- JEQ @SetMem
tmp(177) := "0001" & "000" & "000001011" ;	-- LDA R0, @MEM0
tmp(178) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(179) := "0001" & "001" & "000001100" ;	-- LDA R1, @MEM1
tmp(180) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(181) := "0001" & "010" & "000001101" ;	-- LDA R2, @MEM2
tmp(182) := "0110" & "010" & "100100010" ;	-- STA @HEX2, R2
tmp(183) := "0001" & "011" & "000001110" ;	-- LDA R3, @MEM3
tmp(184) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(185) := "0001" & "111" & "000010001" ;	-- LDA R7, @AMPM
tmp(186) := "1001" & "111" & "000000001" ;	-- CEQ R7, @1
tmp(187) := "1100" & "000" & "010111110" ;	-- JNE @CheckBase24
tmp(188) := "1010" & "000" & "001101110" ;	-- JSR @Base12
tmp(189) := "0111" & "000" & "010111111" ;	-- JMP @KeepWaiting

-- LABEL CheckBase24
tmp(190) := "1010" & "000" & "010001011" ;	-- JSR @Base24

-- LABEL KeepWaiting
tmp(191) := "0001" & "111" & "101100010" ;	-- LDA R7, @KEY2
tmp(192) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(193) := "1001" & "111" & "000000001" ;	-- CEQ R7, @1
tmp(194) := "1100" & "000" & "000111000" ;	-- JNE @IncClk
tmp(195) := "0110" & "000" & "111111101" ;	-- CLR @KEY2
tmp(196) := "0001" & "111" & "000010001" ;	-- LDA R7, @AMPM
tmp(197) := "1001" & "111" & "000000001" ;	-- CEQ R7, @1
tmp(198) := "1000" & "000" & "011001001" ;	-- JEQ @Toggle
tmp(199) := "0001" & "111" & "000000001" ;	-- LDA R7, @1
tmp(200) := "0111" & "000" & "011001010" ;	-- JMP @RetToggle

-- LABEL Toggle
tmp(201) := "0001" & "111" & "000000000" ;	-- LDA R7, @0

-- LABEL RetToggle
tmp(202) := "0110" & "111" & "000010001" ;	-- STA @AMPM, R7
tmp(203) := "0111" & "000" & "000111000" ;	-- JMP @IncClk

-- LABEL SetMem
tmp(204) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(205) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(206) := "0110" & "111" & "100000010" ;	-- STA @LED9, R7
tmp(207) := "0001" & "011" & "000001011" ;	-- LDA R3, @MEM0
tmp(208) := "0110" & "011" & "100100000" ;	-- STA @HEX0, R3
tmp(209) := "0001" & "011" & "000001100" ;	-- LDA R3, @MEM1
tmp(210) := "0110" & "011" & "100100001" ;	-- STA @HEX1, R3
tmp(211) := "0001" & "011" & "000001101" ;	-- LDA R3, @MEM2
tmp(212) := "0110" & "011" & "100100010" ;	-- STA @HEX2, R3
tmp(213) := "0001" & "011" & "000001110" ;	-- LDA R3, @MEM3
tmp(214) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(215) := "0001" & "011" & "000001111" ;	-- LDA R3, @MEM4
tmp(216) := "1110" & "011" & "000000100" ;	-- CLT R3, @4
tmp(217) := "1101" & "000" & "011011100" ;	-- JLT @StartSet4
tmp(218) := "1010" & "000" & "010011000" ;	-- JSR @BAS5SET2
tmp(219) := "0111" & "000" & "011011101" ;	-- JMP @Display4

-- LABEL StartSet4
tmp(220) := "1010" & "000" & "010011011" ;	-- JSR @BAS5SET3

-- LABEL Display4
tmp(221) := "0110" & "011" & "100100100" ;	-- STA @HEX4, R3
tmp(222) := "0001" & "011" & "000010000" ;	-- LDA R3, @MEM5
tmp(223) := "0110" & "011" & "100100101" ;	-- STA @HEX5, R3
tmp(224) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(225) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(226) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(227) := "0001" & "010" & "000000001" ;	-- LDA R2, @1
tmp(228) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(229) := "0110" & "000" & "111111111" ;	-- CLR @KEY0
tmp(230) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(231) := "0111" & "000" & "011101000" ;	-- JMP @VerificaK0

-- LABEL VerificaK0
tmp(232) := "0001" & "110" & "101100000" ;	-- LDA R6, @KEY0
tmp(233) := "0100" & "110" & "000000001" ;	-- AND R6, @1
tmp(234) := "1001" & "110" & "000000000" ;	-- CEQ R6, @0
tmp(235) := "1000" & "000" & "011101101" ;	-- JEQ @VerificaK1
tmp(236) := "0111" & "000" & "011110010" ;	-- JMP @IncMem

-- LABEL VerificaK1
tmp(237) := "0001" & "111" & "101100011" ;	-- LDA R7, @KEY3
tmp(238) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(239) := "1001" & "111" & "000000000" ;	-- CEQ R7, @0
tmp(240) := "1100" & "000" & "100111000" ;	-- JNE @Set0
tmp(241) := "0111" & "000" & "011101000" ;	-- JMP @VerificaK0

-- LABEL IncMem
tmp(242) := "0110" & "000" & "111111111" ;	-- CLR @KEY0
tmp(243) := "1001" & "000" & "000000000" ;	-- CEQ R0, @0
tmp(244) := "1000" & "000" & "011111111" ;	-- JEQ @IncMem0
tmp(245) := "1001" & "000" & "000000001" ;	-- CEQ R0, @1
tmp(246) := "1000" & "000" & "100000111" ;	-- JEQ @IncMem1
tmp(247) := "1001" & "000" & "000000010" ;	-- CEQ R0, @2
tmp(248) := "1000" & "000" & "100001111" ;	-- JEQ @IncMem2
tmp(249) := "1001" & "000" & "000000011" ;	-- CEQ R0, @3
tmp(250) := "1000" & "000" & "100010111" ;	-- JEQ @IncMem3
tmp(251) := "1001" & "000" & "000000100" ;	-- CEQ R0, @4
tmp(252) := "1000" & "000" & "100011111" ;	-- JEQ @IncMem4
tmp(253) := "1001" & "000" & "000000101" ;	-- CEQ R0, @5
tmp(254) := "1000" & "000" & "100101100" ;	-- JEQ @IncMem5

-- LABEL IncMem0
tmp(255) := "0001" & "001" & "000001011" ;	-- LDA R1, @MEM0
tmp(256) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(257) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(258) := "1100" & "000" & "100000100" ;	-- JNE @StaMem0
tmp(259) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem0
tmp(260) := "0110" & "001" & "000001011" ;	-- STA @MEM0, R1
tmp(261) := "0110" & "001" & "100100000" ;	-- STA @HEX0, R1
tmp(262) := "0111" & "000" & "011101101" ;	-- JMP @VerificaK1

-- LABEL IncMem1
tmp(263) := "0001" & "001" & "000001100" ;	-- LDA R1, @MEM1
tmp(264) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(265) := "1001" & "001" & "000000110" ;	-- CEQ R1, @6
tmp(266) := "1100" & "000" & "100001100" ;	-- JNE @StaMem1
tmp(267) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem1
tmp(268) := "0110" & "001" & "000001100" ;	-- STA @MEM1, R1
tmp(269) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(270) := "0111" & "000" & "011101101" ;	-- JMP @VerificaK1

-- LABEL IncMem2
tmp(271) := "0001" & "001" & "000001101" ;	-- LDA R1, @MEM2
tmp(272) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(273) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(274) := "1100" & "000" & "100010100" ;	-- JNE @StaMem2
tmp(275) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem2
tmp(276) := "0110" & "001" & "000001101" ;	-- STA @MEM2, R1
tmp(277) := "0110" & "001" & "100100010" ;	-- STA @HEX2, R1
tmp(278) := "0111" & "000" & "011101101" ;	-- JMP @VerificaK1

-- LABEL IncMem3
tmp(279) := "0001" & "001" & "000001110" ;	-- LDA R1, @MEM3
tmp(280) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(281) := "1001" & "001" & "000000110" ;	-- CEQ R1, @6
tmp(282) := "1100" & "000" & "100011100" ;	-- JNE @StaMem3
tmp(283) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem3
tmp(284) := "0110" & "001" & "000001110" ;	-- STA @MEM3, R1
tmp(285) := "0110" & "001" & "100100011" ;	-- STA @HEX3, R1
tmp(286) := "0111" & "000" & "011101101" ;	-- JMP @VerificaK1

-- LABEL IncMem4
tmp(287) := "0001" & "001" & "000001111" ;	-- LDA R1, @MEM4
tmp(288) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(289) := "1001" & "001" & "000010010" ;	-- CEQ R1, @BAS4
tmp(290) := "1100" & "000" & "100100100" ;	-- JNE @StaMem4
tmp(291) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem4
tmp(292) := "0110" & "001" & "000001111" ;	-- STA @MEM4, R1
tmp(293) := "0110" & "001" & "100100100" ;	-- STA @HEX4, R1
tmp(294) := "1110" & "001" & "000000100" ;	-- CLT R1, @4
tmp(295) := "1101" & "000" & "100101010" ;	-- JLT @setMax3
tmp(296) := "1010" & "000" & "010011000" ;	-- JSR @BAS5SET2
tmp(297) := "0111" & "000" & "011101101" ;	-- JMP @VerificaK1

-- LABEL setMax3
tmp(298) := "1010" & "000" & "010011011" ;	-- JSR @BAS5SET3
tmp(299) := "0111" & "000" & "011101101" ;	-- JMP @VerificaK1

-- LABEL IncMem5
tmp(300) := "0001" & "001" & "000010000" ;	-- LDA R1, @MEM5
tmp(301) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(302) := "1001" & "001" & "000010011" ;	-- CEQ R1, @BAS5
tmp(303) := "1100" & "000" & "100110010" ;	-- JNE @StaMem5
tmp(304) := "0001" & "001" & "000000000" ;	-- LDA R1, $0
tmp(305) := "1010" & "000" & "010010101" ;	-- JSR @BAS4SET10

-- LABEL StaMem5
tmp(306) := "1001" & "001" & "000000010" ;	-- CEQ R1, @2
tmp(307) := "1100" & "000" & "100110101" ;	-- JNE @SetBase24
tmp(308) := "1010" & "000" & "010010010" ;	-- JSR @BAS4SET4

-- LABEL SetBase24
tmp(309) := "0110" & "001" & "000010000" ;	-- STA @MEM5, R1
tmp(310) := "0110" & "001" & "100100101" ;	-- STA @HEX5, R1
tmp(311) := "0111" & "000" & "011101101" ;	-- JMP @VerificaK1

-- LABEL Set0
tmp(312) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(313) := "1001" & "000" & "000000000" ;	-- CEQ R0, @0
tmp(314) := "1000" & "000" & "101010010" ;	-- JEQ @Set1
tmp(315) := "1001" & "000" & "000000001" ;	-- CEQ R0, @1
tmp(316) := "1000" & "000" & "101010110" ;	-- JEQ @Set2
tmp(317) := "1001" & "000" & "000000010" ;	-- CEQ R0, @2
tmp(318) := "1000" & "000" & "101011010" ;	-- JEQ @Set3
tmp(319) := "1001" & "000" & "000000011" ;	-- CEQ R0, @3
tmp(320) := "1000" & "000" & "101011110" ;	-- JEQ @Set4
tmp(321) := "1001" & "000" & "000000100" ;	-- CEQ R0, @4
tmp(322) := "1000" & "000" & "101100010" ;	-- JEQ @Set5
tmp(323) := "0101" & "010" & "000000000" ;	-- LDI R2, @0
tmp(324) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(325) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(326) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(327) := "0001" & "101" & "000000000" ;	-- LDA R5, @0
tmp(328) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(329) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(330) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(331) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(332) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(333) := "0110" & "000" & "111111111" ;	-- CLR @KEY0
tmp(334) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(335) := "0110" & "000" & "111111010" ;	-- CLR @SEC
tmp(336) := "1010" & "000" & "010011011" ;	-- JSR @BAS5SET3
tmp(337) := "0111" & "000" & "000101011" ;	-- JMP @Clock

-- LABEL Set1
tmp(338) := "0101" & "010" & "000000010" ;	-- LDI R2, $2
tmp(339) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(340) := "0101" & "000" & "000000001" ;	-- LDI R0, @1
tmp(341) := "0111" & "000" & "011101000" ;	-- JMP @VerificaK0

-- LABEL Set2
tmp(342) := "0101" & "010" & "000000100" ;	-- LDI R2, $4
tmp(343) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(344) := "0101" & "000" & "000000010" ;	-- LDI R0, @2
tmp(345) := "0111" & "000" & "011101000" ;	-- JMP @VerificaK0

-- LABEL Set3
tmp(346) := "0101" & "010" & "000001000" ;	-- LDI R2, $8
tmp(347) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(348) := "0101" & "000" & "000000011" ;	-- LDI R0, @3
tmp(349) := "0111" & "000" & "011101000" ;	-- JMP @VerificaK0

-- LABEL Set4
tmp(350) := "0101" & "010" & "000010000" ;	-- LDI R2, $16
tmp(351) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(352) := "0101" & "000" & "000000100" ;	-- LDI R0, @4
tmp(353) := "0111" & "000" & "011101000" ;	-- JMP @VerificaK0

-- LABEL Set5
tmp(354) := "0101" & "010" & "000100000" ;	-- LDI R2, $32
tmp(355) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(356) := "0101" & "000" & "000000101" ;	-- LDI R0, @5
tmp(357) := "0111" & "000" & "011101000" ;	-- JMP @VerificaK0

		  
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;