library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 16;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant ANDD : std_logic_vector(3 downto 0) := "0100";
  constant LDI  : std_logic_vector(3 downto 0) := "0101";
  constant STA  : std_logic_vector(3 downto 0) := "0110";
  constant JMP  : std_logic_vector(3 downto 0) := "0111";
  constant JEQ  : std_logic_vector(3 downto 0) := "1000";
  constant CEQ  : std_logic_vector(3 downto 0) := "1001";
  constant JSR  : std_logic_vector(3 downto 0) := "1010";
  constant RET  : std_logic_vector(3 downto 0) := "1011";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
  

-- LABEL Setup
tmp(0) := "0101" & "000" & "000000000" ;	-- LDI R0, $0
tmp(1) := "0110" & "000" & "000000000" ;	-- STA @0, R0
tmp(2) := "0101" & "001" & "000000001" ;	-- LDI R1, $1
tmp(3) := "0110" & "001" & "000000001" ;	-- STA @1, R1
tmp(4) := "0101" & "001" & "000000010" ;	-- LDI R1, $2
tmp(5) := "0110" & "001" & "000000010" ;	-- STA @2, R1
tmp(6) := "0101" & "001" & "000000011" ;	-- LDI R1, $3
tmp(7) := "0110" & "001" & "000000011" ;	-- STA @3, R1
tmp(8) := "0101" & "001" & "000000100" ;	-- LDI R1, $4
tmp(9) := "0110" & "001" & "000000100" ;	-- STA @4, R1
tmp(10) := "0101" & "001" & "000000101" ;	-- LDI R1, $5
tmp(11) := "0110" & "001" & "000000101" ;	-- STA @5, R1
tmp(12) := "0101" & "001" & "000001010" ;	-- LDI R1, $10
tmp(13) := "0110" & "001" & "000001010" ;	-- STA @10, R1
tmp(14) := "0101" & "001" & "000001001" ;	-- LDI R1, $9
tmp(15) := "0110" & "000" & "000010111" ;	-- STA @FLAG, R0
tmp(16) := "0110" & "001" & "000001011" ;	-- STA @LIM0, R1
tmp(17) := "0110" & "001" & "000001100" ;	-- STA @LIM1, R1
tmp(18) := "0110" & "001" & "000001101" ;	-- STA @LIM2, R1
tmp(19) := "0110" & "001" & "000001110" ;	-- STA @LIM3, R1
tmp(20) := "0110" & "001" & "000001111" ;	-- STA @LIM4, R1
tmp(21) := "0110" & "001" & "000010000" ;	-- STA @LIM5, R1
tmp(22) := "0110" & "000" & "000010001" ;	-- STA @MEM0, R0
tmp(23) := "0101" & "001" & "000001000" ;	-- LDI R1, $8
tmp(24) := "0110" & "001" & "000010010" ;	-- STA @MEM1, R1
tmp(25) := "0101" & "001" & "000001001" ;	-- LDI R1, $9
tmp(26) := "0110" & "001" & "000010011" ;	-- STA @MEM2, R1
tmp(27) := "0110" & "000" & "000010100" ;	-- STA @MEM3, R0
tmp(28) := "0110" & "000" & "000010101" ;	-- STA @MEM4, R0
tmp(29) := "0110" & "000" & "000010110" ;	-- STA @MEM5, R0
tmp(30) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(31) := "0110" & "000" & "100100001" ;	-- STA @HEX1, R0
tmp(32) := "0110" & "000" & "100100010" ;	-- STA @HEX2, R0
tmp(33) := "0110" & "000" & "100100011" ;	-- STA @HEX3, R0
tmp(34) := "0110" & "000" & "100100100" ;	-- STA @HEX4, R0
tmp(35) := "0110" & "000" & "100100101" ;	-- STA @HEX5, R0
tmp(36) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(37) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(38) := "0001" & "101" & "000000000" ;	-- LDA R5, @0
tmp(39) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(40) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(41) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(42) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(43) := "0001" & "000" & "000000000" ;	-- LDA R0, @0

-- LABEL Contador
tmp(44) := "0001" & "011" & "000010001" ;	-- LDA R3, @MEM0
tmp(45) := "0110" & "011" & "100100000" ;	-- STA @HEX0, R3
tmp(46) := "0001" & "011" & "000010010" ;	-- LDA R3, @MEM1
tmp(47) := "0110" & "011" & "100100001" ;	-- STA @HEX1, R3
tmp(48) := "0001" & "011" & "000010011" ;	-- LDA R3, @MEM2
tmp(49) := "0110" & "011" & "100100010" ;	-- STA @HEX2, R3
tmp(50) := "0001" & "011" & "000010100" ;	-- LDA R3, @MEM3
tmp(51) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(52) := "0001" & "011" & "000010101" ;	-- LDA R3, @MEM4
tmp(53) := "0110" & "011" & "100100100" ;	-- STA @HEX4, R3
tmp(54) := "0001" & "011" & "000010110" ;	-- LDA R3, @MEM5
tmp(55) := "0110" & "011" & "100100101" ;	-- STA @HEX5, R3
tmp(56) := "0111" & "000" & "000111001" ;	-- JMP @IncCont

-- LABEL IncCont
tmp(57) := "0001" & "110" & "101100010" ;	-- LDA R6, @KEY2
tmp(58) := "0100" & "110" & "000000001" ;	-- AND R6, @1
tmp(59) := "1001" & "110" & "000000001" ;	-- CEQ R6, @1
tmp(60) := "1000" & "000" & "000111110" ;	-- JEQ @IncMem0
tmp(61) := "0111" & "000" & "001110110" ;	-- JMP @WaitLimit

-- LABEL IncMem0
tmp(62) := "0110" & "000" & "111111101" ;	-- CLR @KEY2
tmp(63) := "0001" & "000" & "000010001" ;	-- LDA R0, @MEM0
tmp(64) := "0010" & "000" & "000000001" ;	-- SOMA R0, @1
tmp(65) := "1001" & "000" & "000001010" ;	-- CEQ R0, @10
tmp(66) := "1000" & "000" & "001000110" ;	-- JEQ @ResetMem0
tmp(67) := "0110" & "000" & "000010001" ;	-- STA @MEM0, R0
tmp(68) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(69) := "0111" & "000" & "001111011" ;	-- JMP @Limits

-- LABEL ResetMem0
tmp(70) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(71) := "0110" & "000" & "000010001" ;	-- STA @MEM0, R0
tmp(72) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(73) := "0001" & "001" & "000010010" ;	-- LDA R1, @MEM1
tmp(74) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(75) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(76) := "1000" & "000" & "001010000" ;	-- JEQ @ResetMem1
tmp(77) := "0110" & "001" & "000010010" ;	-- STA @MEM1, R1
tmp(78) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(79) := "0111" & "000" & "001111011" ;	-- JMP @Limits

-- LABEL ResetMem1
tmp(80) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(81) := "0110" & "001" & "000010010" ;	-- STA @MEM1, R1
tmp(82) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(83) := "0001" & "010" & "000010011" ;	-- LDA R2, @MEM2
tmp(84) := "0010" & "010" & "000000001" ;	-- SOMA R2, @1
tmp(85) := "1001" & "010" & "000001010" ;	-- CEQ R2, @10
tmp(86) := "1000" & "000" & "001011010" ;	-- JEQ @ResetMem2
tmp(87) := "0110" & "010" & "000010011" ;	-- STA @MEM2, R2
tmp(88) := "0110" & "010" & "100100010" ;	-- STA @HEX2, R2
tmp(89) := "0111" & "000" & "001111011" ;	-- JMP @Limits

-- LABEL ResetMem2
tmp(90) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(91) := "0110" & "010" & "000010011" ;	-- STA @MEM2, R2
tmp(92) := "0110" & "010" & "100100010" ;	-- STA @HEX2, R2
tmp(93) := "0001" & "011" & "000010100" ;	-- LDA R3, @MEM3
tmp(94) := "0010" & "011" & "000000001" ;	-- SOMA R3, @1
tmp(95) := "1001" & "011" & "000001010" ;	-- CEQ R3, @10
tmp(96) := "1000" & "000" & "001100100" ;	-- JEQ @ResetMem3
tmp(97) := "0110" & "011" & "000010100" ;	-- STA @MEM3, R3
tmp(98) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(99) := "0111" & "000" & "001111011" ;	-- JMP @Limits

-- LABEL ResetMem3
tmp(100) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(101) := "0110" & "011" & "000010100" ;	-- STA @MEM3, R3
tmp(102) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(103) := "0001" & "100" & "000010101" ;	-- LDA R4, @MEM4
tmp(104) := "0010" & "100" & "000000001" ;	-- SOMA R4, @1
tmp(105) := "1001" & "100" & "000001010" ;	-- CEQ R4, @10
tmp(106) := "1000" & "000" & "001101110" ;	-- JEQ @ResetMem4
tmp(107) := "0110" & "100" & "000010101" ;	-- STA @MEM4, R4
tmp(108) := "0110" & "100" & "100100100" ;	-- STA @HEX4, R4
tmp(109) := "0111" & "000" & "001111011" ;	-- JMP @Limits

-- LABEL ResetMem4
tmp(110) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(111) := "0110" & "100" & "000010101" ;	-- STA @MEM4, R4
tmp(112) := "0110" & "100" & "100100100" ;	-- STA @HEX4, R4
tmp(113) := "0001" & "101" & "000010110" ;	-- LDA R5, @MEM5
tmp(114) := "0010" & "101" & "000000001" ;	-- SOMA R5, @1
tmp(115) := "0110" & "101" & "000010110" ;	-- STA @MEM5, R5
tmp(116) := "0110" & "101" & "100100101" ;	-- STA @HEX5, R5
tmp(117) := "0111" & "000" & "001111011" ;	-- JMP @Limits

-- LABEL WaitLimit
tmp(118) := "0001" & "111" & "101100011" ;	-- LDA R7, @KEY3
tmp(119) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(120) := "1001" & "111" & "000000001" ;	-- CEQ R7, @1
tmp(121) := "1000" & "000" & "010101111" ;	-- JEQ @SetLimit
tmp(122) := "0111" & "000" & "000111001" ;	-- JMP @IncCont

-- LABEL Limits
tmp(123) := "1010" & "000" & "001111110" ;	-- JSR @Limiter5
tmp(124) := "1010" & "000" & "010011011" ;	-- JSR @VerificaFlag
tmp(125) := "0111" & "000" & "001110110" ;	-- JMP @WaitLimit

-- LABEL Limiter5
tmp(126) := "0001" & "000" & "000010000" ;	-- LDA R0, @LIM5
tmp(127) := "1001" & "000" & "000010110" ;	-- CEQ R0, @MEM5
tmp(128) := "1000" & "000" & "010000010" ;	-- JEQ @Limiter4
tmp(129) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Limiter4
tmp(130) := "0001" & "000" & "000001111" ;	-- LDA R0, @LIM4
tmp(131) := "1001" & "000" & "000010101" ;	-- CEQ R0, @MEM4
tmp(132) := "1000" & "000" & "010000110" ;	-- JEQ @Limiter3
tmp(133) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Limiter3
tmp(134) := "0001" & "000" & "000001110" ;	-- LDA R0, @LIM3
tmp(135) := "1001" & "000" & "000010100" ;	-- CEQ R0, @MEM3
tmp(136) := "1000" & "000" & "010001010" ;	-- JEQ @Limiter2
tmp(137) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Limiter2
tmp(138) := "0001" & "000" & "000001101" ;	-- LDA R0, @LIM2
tmp(139) := "1001" & "000" & "000010011" ;	-- CEQ R0, @MEM2
tmp(140) := "1000" & "000" & "010001110" ;	-- JEQ @Limiter1
tmp(141) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Limiter1
tmp(142) := "0001" & "000" & "000001100" ;	-- LDA R0, @LIM1
tmp(143) := "1001" & "000" & "000010010" ;	-- CEQ R0, @MEM1
tmp(144) := "1000" & "000" & "010010010" ;	-- JEQ @Limiter0
tmp(145) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Limiter0
tmp(146) := "0001" & "000" & "000001011" ;	-- LDA R0, @LIM0
tmp(147) := "1001" & "000" & "000010001" ;	-- CEQ R0, @MEM0
tmp(148) := "1000" & "000" & "010010110" ;	-- JEQ @AcionaFlag
tmp(149) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL AcionaFlag
tmp(150) := "0001" & "000" & "000000001" ;	-- LDA R0, @1
tmp(151) := "0110" & "000" & "000010111" ;	-- STA @FLAG, R0
tmp(152) := "0110" & "000" & "100000010" ;	-- STA @LED9, R0
tmp(153) := "0110" & "000" & "100000001" ;	-- STA @LED8, R0
tmp(154) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL VerificaFlag
tmp(155) := "0001" & "000" & "000000001" ;	-- LDA R0, @1
tmp(156) := "1001" & "000" & "000010111" ;	-- CEQ R0, @FLAG
tmp(157) := "1000" & "000" & "010011111" ;	-- JEQ @Parado
tmp(158) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Parado
tmp(159) := "0001" & "000" & "101100011" ;	-- LDA R0, @KEY3
tmp(160) := "0100" & "000" & "000000001" ;	-- AND R0, @1
tmp(161) := "1001" & "000" & "000000001" ;	-- CEQ R0, @1
tmp(162) := "1000" & "000" & "010101111" ;	-- JEQ @SetLimit
tmp(163) := "0001" & "000" & "101100010" ;	-- LDA R0, @KEY2
tmp(164) := "0100" & "000" & "000000001" ;	-- AND R0, @1
tmp(165) := "1001" & "000" & "000000001" ;	-- CEQ R0, @1
tmp(166) := "1000" & "000" & "010101000" ;	-- JEQ @AllLEDs
tmp(167) := "0111" & "000" & "010011111" ;	-- JMP @Parado

-- LABEL AllLEDs
tmp(168) := "0110" & "000" & "111111101" ;	-- CLR @KEY2
tmp(169) := "0101" & "001" & "011111111" ;	-- LDI R1, $255
tmp(170) := "0110" & "001" & "100000000" ;	-- STA @LEDb, R1
tmp(171) := "0101" & "001" & "000000001" ;	-- LDI R1, $1
tmp(172) := "0110" & "001" & "100000001" ;	-- STA @LED8, R1
tmp(173) := "0110" & "001" & "100000010" ;	-- STA @LED9, R1
tmp(174) := "0111" & "000" & "010011111" ;	-- JMP @Parado

-- LABEL SetLimit
tmp(175) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(176) := "0001" & "011" & "000001011" ;	-- LDA R3, @LIM0
tmp(177) := "0110" & "011" & "100100000" ;	-- STA @HEX0, R3
tmp(178) := "0001" & "011" & "000001100" ;	-- LDA R3, @LIM1
tmp(179) := "0110" & "011" & "100100001" ;	-- STA @HEX1, R3
tmp(180) := "0001" & "011" & "000001101" ;	-- LDA R3, @LIM2
tmp(181) := "0110" & "011" & "100100010" ;	-- STA @HEX2, R3
tmp(182) := "0001" & "011" & "000001110" ;	-- LDA R3, @LIM3
tmp(183) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(184) := "0001" & "011" & "000001111" ;	-- LDA R3, @LIM4
tmp(185) := "0110" & "011" & "100100100" ;	-- STA @HEX4, R3
tmp(186) := "0001" & "011" & "000010000" ;	-- LDA R3, @LIM5
tmp(187) := "0110" & "011" & "100100101" ;	-- STA @HEX5, R3
tmp(188) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(189) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(190) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(191) := "0110" & "000" & "100000001" ;	-- STA @LED8, R0
tmp(192) := "0110" & "000" & "100000010" ;	-- STA @LED9, R0
tmp(193) := "0001" & "010" & "000000001" ;	-- LDA R2, @1
tmp(194) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(195) := "0110" & "000" & "111111111" ;	-- CLR @KEY0
tmp(196) := "0110" & "000" & "111111110" ;	-- CLR @KEY1
tmp(197) := "0111" & "000" & "011000110" ;	-- JMP @VerificaK0

-- LABEL VerificaK0
tmp(198) := "0001" & "110" & "101100000" ;	-- LDA R6, @KEY0
tmp(199) := "0100" & "110" & "000000001" ;	-- AND R6, @1
tmp(200) := "1001" & "110" & "000000000" ;	-- CEQ R6, @0
tmp(201) := "1000" & "000" & "011001011" ;	-- JEQ @VerificaK1
tmp(202) := "1010" & "000" & "011010001" ;	-- JSR @IncLim

-- LABEL VerificaK1
tmp(203) := "0001" & "111" & "101100001" ;	-- LDA R7, @KEY1
tmp(204) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(205) := "1001" & "111" & "000000000" ;	-- CEQ R7, @0
tmp(206) := "1000" & "000" & "011000110" ;	-- JEQ @VerificaK0
tmp(207) := "1010" & "000" & "100010100" ;	-- JSR @Set0
tmp(208) := "0111" & "000" & "011000110" ;	-- JMP @VerificaK0

-- LABEL IncLim
tmp(209) := "0110" & "000" & "111111111" ;	-- CLR @KEY0
tmp(210) := "1001" & "000" & "000000000" ;	-- CEQ R0, @0
tmp(211) := "1000" & "000" & "011011110" ;	-- JEQ @IncLim0
tmp(212) := "1001" & "000" & "000000001" ;	-- CEQ R0, @1
tmp(213) := "1000" & "000" & "011100111" ;	-- JEQ @IncLim1
tmp(214) := "1001" & "000" & "000000010" ;	-- CEQ R0, @2
tmp(215) := "1000" & "000" & "011110000" ;	-- JEQ @IncLim2
tmp(216) := "1001" & "000" & "000000011" ;	-- CEQ R0, @3
tmp(217) := "1000" & "000" & "011111001" ;	-- JEQ @IncLim3
tmp(218) := "1001" & "000" & "000000100" ;	-- CEQ R0, @4
tmp(219) := "1000" & "000" & "100000010" ;	-- JEQ @IncLim4
tmp(220) := "1001" & "000" & "000000101" ;	-- CEQ R0, @5
tmp(221) := "1000" & "000" & "100001011" ;	-- JEQ @IncLim5

-- LABEL IncLim0
tmp(222) := "0001" & "001" & "000001011" ;	-- LDA R1, @LIM0
tmp(223) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(224) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(225) := "1000" & "000" & "011100011" ;	-- JEQ @ResetLim0
tmp(226) := "0111" & "000" & "011100100" ;	-- JMP @StaLim0

-- LABEL ResetLim0
tmp(227) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaLim0
tmp(228) := "0110" & "001" & "000001011" ;	-- STA @LIM0, R1
tmp(229) := "0110" & "001" & "100100000" ;	-- STA @HEX0, R1
tmp(230) := "0111" & "000" & "011001011" ;	-- JMP @VerificaK1

-- LABEL IncLim1
tmp(231) := "0001" & "001" & "000001100" ;	-- LDA R1, @LIM1
tmp(232) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(233) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(234) := "1000" & "000" & "011101100" ;	-- JEQ @ResetLim1
tmp(235) := "0111" & "000" & "011101101" ;	-- JMP @StaLim1

-- LABEL ResetLim1
tmp(236) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaLim1
tmp(237) := "0110" & "001" & "000001100" ;	-- STA @LIM1, R1
tmp(238) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(239) := "0111" & "000" & "011001011" ;	-- JMP @VerificaK1

-- LABEL IncLim2
tmp(240) := "0001" & "001" & "000001101" ;	-- LDA R1, @LIM2
tmp(241) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(242) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(243) := "1000" & "000" & "011110101" ;	-- JEQ @ResetLim2
tmp(244) := "0111" & "000" & "011110110" ;	-- JMP @StaLim2

-- LABEL ResetLim2
tmp(245) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaLim2
tmp(246) := "0110" & "001" & "000001101" ;	-- STA @LIM2, R1
tmp(247) := "0110" & "001" & "100100010" ;	-- STA @HEX2, R1
tmp(248) := "0111" & "000" & "011001011" ;	-- JMP @VerificaK1

-- LABEL IncLim3
tmp(249) := "0001" & "001" & "000001110" ;	-- LDA R1, @LIM3
tmp(250) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(251) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(252) := "1000" & "000" & "011111110" ;	-- JEQ @ResetLim3
tmp(253) := "0111" & "000" & "011111111" ;	-- JMP @StaLim3

-- LABEL ResetLim3
tmp(254) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaLim3
tmp(255) := "0110" & "001" & "000001110" ;	-- STA @LIM3, R1
tmp(256) := "0110" & "001" & "100100011" ;	-- STA @HEX3, R1
tmp(257) := "0111" & "000" & "011001011" ;	-- JMP @VerificaK1

-- LABEL IncLim4
tmp(258) := "0001" & "001" & "000001111" ;	-- LDA R1, @LIM4
tmp(259) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(260) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(261) := "1000" & "000" & "100000111" ;	-- JEQ @ResetLim4
tmp(262) := "0111" & "000" & "100001000" ;	-- JMP @StaLim4

-- LABEL ResetLim4
tmp(263) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaLim4
tmp(264) := "0110" & "001" & "000001111" ;	-- STA @LIM4, R1
tmp(265) := "0110" & "001" & "100100100" ;	-- STA @HEX4, R1
tmp(266) := "0111" & "000" & "011001011" ;	-- JMP @VerificaK1

-- LABEL IncLim5
tmp(267) := "0001" & "001" & "000010000" ;	-- LDA R1, @LIM5
tmp(268) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(269) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(270) := "1000" & "000" & "100010000" ;	-- JEQ @ResetLim5
tmp(271) := "0111" & "000" & "100010001" ;	-- JMP @StaLim5

-- LABEL ResetLim5
tmp(272) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaLim5
tmp(273) := "0110" & "001" & "000010000" ;	-- STA @LIM5, R1
tmp(274) := "0110" & "001" & "100100101" ;	-- STA @HEX5, R1
tmp(275) := "0111" & "000" & "011001011" ;	-- JMP @VerificaK1

-- LABEL Set0
tmp(276) := "0110" & "000" & "111111110" ;	-- CLR @KEY1
tmp(277) := "1001" & "000" & "000000000" ;	-- CEQ R0, @0
tmp(278) := "1000" & "000" & "100101101" ;	-- JEQ @Set1
tmp(279) := "1001" & "000" & "000000001" ;	-- CEQ R0, @1
tmp(280) := "1000" & "000" & "100110001" ;	-- JEQ @Set2
tmp(281) := "1001" & "000" & "000000010" ;	-- CEQ R0, @2
tmp(282) := "1000" & "000" & "100110101" ;	-- JEQ @Set3
tmp(283) := "1001" & "000" & "000000011" ;	-- CEQ R0, @3
tmp(284) := "1000" & "000" & "100111001" ;	-- JEQ @Set4
tmp(285) := "1001" & "000" & "000000100" ;	-- CEQ R0, @4
tmp(286) := "1000" & "000" & "100111101" ;	-- JEQ @Set5
tmp(287) := "0101" & "010" & "000000000" ;	-- LDI R2, @0
tmp(288) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(289) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(290) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(291) := "0001" & "101" & "000000000" ;	-- LDA R5, @0
tmp(292) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(293) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(294) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(295) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(296) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(297) := "0110" & "000" & "111111101" ;	-- CLR @KEY2
tmp(298) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(299) := "0110" & "000" & "000010111" ;	-- STA @FLAG, R0
tmp(300) := "0111" & "000" & "000101100" ;	-- JMP @Contador

-- LABEL Set1
tmp(301) := "0101" & "010" & "000000010" ;	-- LDI R2, $2
tmp(302) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(303) := "0101" & "000" & "000000001" ;	-- LDI R0, @1
tmp(304) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Set2
tmp(305) := "0101" & "010" & "000000100" ;	-- LDI R2, $4
tmp(306) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(307) := "0101" & "000" & "000000010" ;	-- LDI R0, @2
tmp(308) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Set3
tmp(309) := "0101" & "010" & "000001000" ;	-- LDI R2, $8
tmp(310) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(311) := "0101" & "000" & "000000011" ;	-- LDI R0, @3
tmp(312) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Set4
tmp(313) := "0101" & "010" & "000010000" ;	-- LDI R2, $16
tmp(314) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(315) := "0101" & "000" & "000000100" ;	-- LDI R0, @4
tmp(316) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Set5
tmp(317) := "0101" & "010" & "000100000" ;	-- LDI R2, $32
tmp(318) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(319) := "0101" & "000" & "000000101" ;	-- LDI R0, @5
tmp(320) := "1011" & "000" & "000000000" ;	-- RET

		  
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;