library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 16;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant ANDD : std_logic_vector(3 downto 0) := "0100";
  constant LDI  : std_logic_vector(3 downto 0) := "0101";
  constant STA  : std_logic_vector(3 downto 0) := "0110";
  constant JMP  : std_logic_vector(3 downto 0) := "0111";
  constant JEQ  : std_logic_vector(3 downto 0) := "1000";
  constant CEQ  : std_logic_vector(3 downto 0) := "1001";
  constant JSR  : std_logic_vector(3 downto 0) := "1010";
  constant RET  : std_logic_vector(3 downto 0) := "1011";
  constant JNE  : std_logic_vector(3 downto 0) := "1100";
  constant JLT  : std_logic_vector(3 downto 0) := "1101";
  constant CLT  : std_logic_vector(3 downto 0) := "1110";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
  

-- LABEL Setup
tmp(0) := "0101" & "000" & "010000000" ;	-- LDI R0, $128
tmp(1) := "0110" & "000" & "000111111" ;	-- STA @63, R0
tmp(2) := "0101" & "000" & "000000000" ;	-- LDI R0, $0
tmp(3) := "0110" & "000" & "000000000" ;	-- STA @0, R0
tmp(4) := "0101" & "001" & "000000001" ;	-- LDI R1, $1
tmp(5) := "0110" & "001" & "000000001" ;	-- STA @1, R1
tmp(6) := "0101" & "001" & "000000010" ;	-- LDI R1, $2
tmp(7) := "0110" & "001" & "000000010" ;	-- STA @2, R1
tmp(8) := "0101" & "001" & "000000011" ;	-- LDI R1, $3
tmp(9) := "0110" & "001" & "000000011" ;	-- STA @3, R1
tmp(10) := "0110" & "001" & "000011001" ;	-- STA @BAS5, R1
tmp(11) := "0101" & "001" & "000000100" ;	-- LDI R1, $4
tmp(12) := "0110" & "001" & "000000100" ;	-- STA @4, R1
tmp(13) := "0101" & "001" & "000000101" ;	-- LDI R1, $5
tmp(14) := "0110" & "001" & "000000101" ;	-- STA @5, R1
tmp(15) := "0101" & "001" & "000000110" ;	-- LDI R1, $6
tmp(16) := "0110" & "001" & "000000110" ;	-- STA @6, R1
tmp(17) := "0101" & "001" & "000001010" ;	-- LDI R1, $10
tmp(18) := "0110" & "001" & "000001010" ;	-- STA @10, R1
tmp(19) := "0110" & "001" & "000011000" ;	-- STA @BAS4, R1
tmp(20) := "0101" & "001" & "000001001" ;	-- LDI R1, $9
tmp(21) := "0110" & "000" & "000010001" ;	-- STA @MEM0, R0
tmp(22) := "0110" & "000" & "000010011" ;	-- STA @MEM2, R0
tmp(23) := "0110" & "000" & "000010010" ;	-- STA @MEM1, R0
tmp(24) := "0110" & "000" & "000010100" ;	-- STA @MEM3, R0
tmp(25) := "0110" & "000" & "000010101" ;	-- STA @MEM4, R0
tmp(26) := "0110" & "000" & "000010110" ;	-- STA @MEM5, R0
tmp(27) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(28) := "0110" & "000" & "100100001" ;	-- STA @HEX1, R0
tmp(29) := "0110" & "000" & "100100010" ;	-- STA @HEX2, R0
tmp(30) := "0110" & "000" & "100100011" ;	-- STA @HEX3, R0
tmp(31) := "0110" & "000" & "100100100" ;	-- STA @HEX4, R0
tmp(32) := "0110" & "000" & "100100101" ;	-- STA @HEX5, R0
tmp(33) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(34) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(35) := "0001" & "101" & "000000000" ;	-- LDA R5, @0
tmp(36) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(37) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(38) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(39) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(40) := "0001" & "000" & "000000000" ;	-- LDA R0, @0

-- LABEL Clock
tmp(41) := "0001" & "011" & "000010001" ;	-- LDA R3, @MEM0
tmp(42) := "0110" & "011" & "100100000" ;	-- STA @HEX0, R3
tmp(43) := "0001" & "011" & "000010010" ;	-- LDA R3, @MEM1
tmp(44) := "0110" & "011" & "100100001" ;	-- STA @HEX1, R3
tmp(45) := "0001" & "011" & "000010011" ;	-- LDA R3, @MEM2
tmp(46) := "0110" & "011" & "100100010" ;	-- STA @HEX2, R3
tmp(47) := "0001" & "011" & "000010100" ;	-- LDA R3, @MEM3
tmp(48) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(49) := "0001" & "011" & "000010101" ;	-- LDA R3, @MEM4
tmp(50) := "0110" & "011" & "100100100" ;	-- STA @HEX4, R3
tmp(51) := "0001" & "011" & "000010110" ;	-- LDA R3, @MEM5
tmp(52) := "0110" & "011" & "100100101" ;	-- STA @HEX5, R3
tmp(53) := "0111" & "000" & "000110110" ;	-- JMP @IncClk

-- LABEL IncClk
tmp(54) := "0001" & "111" & "101100101" ;	-- LDA R7, @SEC
tmp(55) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(56) := "1001" & "111" & "000000001" ;	-- CEQ R7, @1
tmp(57) := "1100" & "000" & "010010001" ;	-- JNE @WaitSet
tmp(58) := "0110" & "000" & "111111010" ;	-- CLR @SEC
tmp(59) := "0001" & "000" & "000010001" ;	-- LDA R0, @MEM0
tmp(60) := "0010" & "000" & "000000001" ;	-- SOMA R0, @1
tmp(61) := "1001" & "000" & "000001010" ;	-- CEQ R0, @10
tmp(62) := "1000" & "000" & "001000010" ;	-- JEQ @ResetMem0
tmp(63) := "0110" & "000" & "000010001" ;	-- STA @MEM0, R0
tmp(64) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(65) := "0111" & "000" & "010010001" ;	-- JMP @WaitSet

-- LABEL ResetMem0
tmp(66) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(67) := "0110" & "000" & "000010001" ;	-- STA @MEM0, R0
tmp(68) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(69) := "0001" & "001" & "000010010" ;	-- LDA R1, @MEM1
tmp(70) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(71) := "1001" & "001" & "000000110" ;	-- CEQ R1, @6
tmp(72) := "1000" & "000" & "001001100" ;	-- JEQ @ResetMem1
tmp(73) := "0110" & "001" & "000010010" ;	-- STA @MEM1, R1
tmp(74) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(75) := "0111" & "000" & "010010001" ;	-- JMP @WaitSet

-- LABEL ResetMem1
tmp(76) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(77) := "0110" & "001" & "000010010" ;	-- STA @MEM1, R1
tmp(78) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(79) := "0001" & "010" & "000010011" ;	-- LDA R2, @MEM2
tmp(80) := "0010" & "010" & "000000001" ;	-- SOMA R2, @1
tmp(81) := "1001" & "010" & "000001010" ;	-- CEQ R2, @10
tmp(82) := "1000" & "000" & "001010110" ;	-- JEQ @ResetMem2
tmp(83) := "0110" & "010" & "000010011" ;	-- STA @MEM2, R2
tmp(84) := "0110" & "010" & "100100010" ;	-- STA @HEX2, R2
tmp(85) := "0111" & "000" & "010010001" ;	-- JMP @WaitSet

-- LABEL ResetMem2
tmp(86) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(87) := "0110" & "010" & "000010011" ;	-- STA @MEM2, R2
tmp(88) := "0110" & "010" & "100100010" ;	-- STA @HEX2, R2
tmp(89) := "0001" & "011" & "000010100" ;	-- LDA R3, @MEM3
tmp(90) := "0010" & "011" & "000000001" ;	-- SOMA R3, @1
tmp(91) := "1001" & "011" & "000000110" ;	-- CEQ R3, @6
tmp(92) := "1000" & "000" & "001100000" ;	-- JEQ @ResetMem3
tmp(93) := "0110" & "011" & "000010100" ;	-- STA @MEM3, R3
tmp(94) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(95) := "0111" & "000" & "010010001" ;	-- JMP @WaitSet

-- LABEL ResetMem3
tmp(96) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(97) := "0110" & "011" & "000010100" ;	-- STA @MEM3, R3
tmp(98) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(99) := "0001" & "100" & "000010101" ;	-- LDA R4, @MEM4
tmp(100) := "0010" & "100" & "000000001" ;	-- SOMA R4, @1
tmp(101) := "1001" & "100" & "000011000" ;	-- CEQ R4, @BAS4
tmp(102) := "1000" & "000" & "001101010" ;	-- JEQ @ResetMem4
tmp(103) := "0110" & "100" & "000010101" ;	-- STA @MEM4, R4
tmp(104) := "0110" & "100" & "100100100" ;	-- STA @HEX4, R4
tmp(105) := "0111" & "000" & "010010001" ;	-- JMP @WaitSet

-- LABEL ResetMem4
tmp(106) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(107) := "0110" & "100" & "000010101" ;	-- STA @MEM4, R4
tmp(108) := "0110" & "100" & "100100100" ;	-- STA @HEX4, R4
tmp(109) := "0001" & "101" & "000010110" ;	-- LDA R5, @MEM5
tmp(110) := "0010" & "101" & "000000001" ;	-- SOMA R5, @1
tmp(111) := "1001" & "101" & "000011001" ;	-- CEQ R5, @BAS5
tmp(112) := "1000" & "000" & "010000010" ;	-- JEQ @Zera
tmp(113) := "0110" & "101" & "000010110" ;	-- STA @MEM5, R5
tmp(114) := "0110" & "101" & "100100101" ;	-- STA @HEX5, R5
tmp(115) := "1001" & "101" & "000000010" ;	-- CEQ R5, @2
tmp(116) := "1010" & "000" & "001110110" ;	-- JSR @BAS4SET4
tmp(117) := "0111" & "000" & "010010001" ;	-- JMP @WaitSet

-- LABEL BAS4SET4
tmp(118) := "0001" & "100" & "000000100" ;	-- LDA R4, @4
tmp(119) := "0110" & "100" & "000011000" ;	-- STA @BAS4, R4
tmp(120) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL BAS4SET10
tmp(121) := "0001" & "100" & "000001010" ;	-- LDA R4, @10
tmp(122) := "0110" & "100" & "000011000" ;	-- STA @BAS4, R4
tmp(123) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL BAS5SET2
tmp(124) := "0001" & "100" & "000000010" ;	-- LDA R4, @2
tmp(125) := "0110" & "100" & "000011001" ;	-- STA @BAS5, R4
tmp(126) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL BAS5SET3
tmp(127) := "0001" & "100" & "000000011" ;	-- LDA R4, @3
tmp(128) := "0110" & "100" & "000011001" ;	-- STA @BAS5, R4
tmp(129) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Zera
tmp(130) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(131) := "0110" & "000" & "000010001" ;	-- STA @MEM0, R0
tmp(132) := "0110" & "000" & "000010011" ;	-- STA @MEM2, R0
tmp(133) := "0110" & "000" & "000010010" ;	-- STA @MEM1, R0
tmp(134) := "0110" & "000" & "000010100" ;	-- STA @MEM3, R0
tmp(135) := "0110" & "000" & "000010101" ;	-- STA @MEM4, R0
tmp(136) := "0110" & "000" & "000010110" ;	-- STA @MEM5, R0
tmp(137) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(138) := "0110" & "000" & "100100001" ;	-- STA @HEX1, R0
tmp(139) := "0110" & "000" & "100100010" ;	-- STA @HEX2, R0
tmp(140) := "0110" & "000" & "100100011" ;	-- STA @HEX3, R0
tmp(141) := "0110" & "000" & "100100100" ;	-- STA @HEX4, R0
tmp(142) := "0110" & "000" & "100100101" ;	-- STA @HEX5, R0
tmp(143) := "1010" & "000" & "001111001" ;	-- JSR @BAS4SET10
tmp(144) := "0111" & "000" & "010010001" ;	-- JMP @WaitSet

-- LABEL WaitSet
tmp(145) := "0001" & "111" & "101100011" ;	-- LDA R7, @KEY3
tmp(146) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(147) := "1001" & "111" & "000000001" ;	-- CEQ R7, @1
tmp(148) := "1000" & "000" & "010010110" ;	-- JEQ @SetMem
tmp(149) := "0111" & "000" & "000110110" ;	-- JMP @IncClk

-- LABEL SetMem
tmp(150) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(151) := "0001" & "011" & "000010001" ;	-- LDA R3, @MEM0
tmp(152) := "0110" & "011" & "100100000" ;	-- STA @HEX0, R3
tmp(153) := "0001" & "011" & "000010010" ;	-- LDA R3, @MEM1
tmp(154) := "0110" & "011" & "100100001" ;	-- STA @HEX1, R3
tmp(155) := "0001" & "011" & "000010011" ;	-- LDA R3, @MEM2
tmp(156) := "0110" & "011" & "100100010" ;	-- STA @HEX2, R3
tmp(157) := "0001" & "011" & "000010100" ;	-- LDA R3, @MEM3
tmp(158) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(159) := "0001" & "011" & "000010101" ;	-- LDA R3, @MEM4
tmp(160) := "1110" & "011" & "000000100" ;	-- CLT R3, @4
tmp(161) := "1101" & "000" & "010100100" ;	-- JLT @StartSet4
tmp(162) := "1010" & "000" & "001111100" ;	-- JSR @BAS5SET2
tmp(163) := "0111" & "000" & "010100101" ;	-- JMP @Display4

-- LABEL StartSet4
tmp(164) := "1010" & "000" & "001111111" ;	-- JSR @BAS5SET3

-- LABEL Display4
tmp(165) := "0110" & "011" & "100100100" ;	-- STA @HEX4, R3
tmp(166) := "0001" & "011" & "000010110" ;	-- LDA R3, @MEM5
tmp(167) := "0110" & "011" & "100100101" ;	-- STA @HEX5, R3
tmp(168) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(169) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(170) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(171) := "0001" & "010" & "000000001" ;	-- LDA R2, @1
tmp(172) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(173) := "0110" & "000" & "111111111" ;	-- CLR @KEY0
tmp(174) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(175) := "0111" & "000" & "010110000" ;	-- JMP @VerificaK0

-- LABEL VerificaK0
tmp(176) := "0001" & "110" & "101100000" ;	-- LDA R6, @KEY0
tmp(177) := "0100" & "110" & "000000001" ;	-- AND R6, @1
tmp(178) := "1001" & "110" & "000000000" ;	-- CEQ R6, @0
tmp(179) := "1000" & "000" & "010110101" ;	-- JEQ @VerificaK1
tmp(180) := "0111" & "000" & "010111010" ;	-- JMP @IncMem

-- LABEL VerificaK1
tmp(181) := "0001" & "111" & "101100011" ;	-- LDA R7, @KEY3
tmp(182) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(183) := "1001" & "111" & "000000000" ;	-- CEQ R7, @0
tmp(184) := "1100" & "000" & "100000000" ;	-- JNE @Set0
tmp(185) := "0111" & "000" & "010110000" ;	-- JMP @VerificaK0

-- LABEL IncMem
tmp(186) := "0110" & "000" & "111111111" ;	-- CLR @KEY0
tmp(187) := "1001" & "000" & "000000000" ;	-- CEQ R0, @0
tmp(188) := "1000" & "000" & "011000111" ;	-- JEQ @IncMem0
tmp(189) := "1001" & "000" & "000000001" ;	-- CEQ R0, @1
tmp(190) := "1000" & "000" & "011001111" ;	-- JEQ @IncMem1
tmp(191) := "1001" & "000" & "000000010" ;	-- CEQ R0, @2
tmp(192) := "1000" & "000" & "011010111" ;	-- JEQ @IncMem2
tmp(193) := "1001" & "000" & "000000011" ;	-- CEQ R0, @3
tmp(194) := "1000" & "000" & "011011111" ;	-- JEQ @IncMem3
tmp(195) := "1001" & "000" & "000000100" ;	-- CEQ R0, @4
tmp(196) := "1000" & "000" & "011100111" ;	-- JEQ @IncMem4
tmp(197) := "1001" & "000" & "000000101" ;	-- CEQ R0, @5
tmp(198) := "1000" & "000" & "011110100" ;	-- JEQ @IncMem5

-- LABEL IncMem0
tmp(199) := "0001" & "001" & "000010001" ;	-- LDA R1, @MEM0
tmp(200) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(201) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(202) := "1100" & "000" & "011001100" ;	-- JNE @StaMem0
tmp(203) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem0
tmp(204) := "0110" & "001" & "000010001" ;	-- STA @MEM0, R1
tmp(205) := "0110" & "001" & "100100000" ;	-- STA @HEX0, R1
tmp(206) := "0111" & "000" & "010110101" ;	-- JMP @VerificaK1

-- LABEL IncMem1
tmp(207) := "0001" & "001" & "000010010" ;	-- LDA R1, @MEM1
tmp(208) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(209) := "1001" & "001" & "000000110" ;	-- CEQ R1, @6
tmp(210) := "1100" & "000" & "011010100" ;	-- JNE @StaMem1
tmp(211) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem1
tmp(212) := "0110" & "001" & "000010010" ;	-- STA @MEM1, R1
tmp(213) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(214) := "0111" & "000" & "010110101" ;	-- JMP @VerificaK1

-- LABEL IncMem2
tmp(215) := "0001" & "001" & "000010011" ;	-- LDA R1, @MEM2
tmp(216) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(217) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(218) := "1100" & "000" & "011011100" ;	-- JNE @StaMem2
tmp(219) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem2
tmp(220) := "0110" & "001" & "000010011" ;	-- STA @MEM2, R1
tmp(221) := "0110" & "001" & "100100010" ;	-- STA @HEX2, R1
tmp(222) := "0111" & "000" & "010110101" ;	-- JMP @VerificaK1

-- LABEL IncMem3
tmp(223) := "0001" & "001" & "000010100" ;	-- LDA R1, @MEM3
tmp(224) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(225) := "1001" & "001" & "000000110" ;	-- CEQ R1, @6
tmp(226) := "1100" & "000" & "011100100" ;	-- JNE @StaMem3
tmp(227) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem3
tmp(228) := "0110" & "001" & "000010100" ;	-- STA @MEM3, R1
tmp(229) := "0110" & "001" & "100100011" ;	-- STA @HEX3, R1
tmp(230) := "0111" & "000" & "010110101" ;	-- JMP @VerificaK1

-- LABEL IncMem4
tmp(231) := "0001" & "001" & "000010101" ;	-- LDA R1, @MEM4
tmp(232) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(233) := "1001" & "001" & "000011000" ;	-- CEQ R1, @BAS4
tmp(234) := "1100" & "000" & "011101100" ;	-- JNE @StaMem4
tmp(235) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem4
tmp(236) := "0110" & "001" & "000010101" ;	-- STA @MEM4, R1
tmp(237) := "0110" & "001" & "100100100" ;	-- STA @HEX4, R1
tmp(238) := "1110" & "001" & "000000100" ;	-- CLT R1, @4
tmp(239) := "1101" & "000" & "011110010" ;	-- JLT @setMax3
tmp(240) := "1010" & "000" & "001111100" ;	-- JSR @BAS5SET2
tmp(241) := "0111" & "000" & "010110101" ;	-- JMP @VerificaK1

-- LABEL setMax3
tmp(242) := "1010" & "000" & "001111111" ;	-- JSR @BAS5SET3
tmp(243) := "0111" & "000" & "010110101" ;	-- JMP @VerificaK1

-- LABEL IncMem5
tmp(244) := "0001" & "001" & "000010110" ;	-- LDA R1, @MEM5
tmp(245) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(246) := "1001" & "001" & "000011001" ;	-- CEQ R1, @BAS5
tmp(247) := "1100" & "000" & "011111010" ;	-- JNE @StaMem5
tmp(248) := "0001" & "001" & "000000000" ;	-- LDA R1, $0
tmp(249) := "1010" & "000" & "001111001" ;	-- JSR @BAS4SET10

-- LABEL StaMem5
tmp(250) := "1001" & "001" & "000000010" ;	-- CEQ R1, @2
tmp(251) := "1100" & "000" & "011111101" ;	-- JNE @SetBase24
tmp(252) := "1010" & "000" & "001110110" ;	-- JSR @BAS4SET4

-- LABEL SetBase24
tmp(253) := "0110" & "001" & "000010110" ;	-- STA @MEM5, R1
tmp(254) := "0110" & "001" & "100100101" ;	-- STA @HEX5, R1
tmp(255) := "0111" & "000" & "010110101" ;	-- JMP @VerificaK1

-- LABEL Set0
tmp(256) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(257) := "1001" & "000" & "000000000" ;	-- CEQ R0, @0
tmp(258) := "1000" & "000" & "100011010" ;	-- JEQ @Set1
tmp(259) := "1001" & "000" & "000000001" ;	-- CEQ R0, @1
tmp(260) := "1000" & "000" & "100011110" ;	-- JEQ @Set2
tmp(261) := "1001" & "000" & "000000010" ;	-- CEQ R0, @2
tmp(262) := "1000" & "000" & "100100010" ;	-- JEQ @Set3
tmp(263) := "1001" & "000" & "000000011" ;	-- CEQ R0, @3
tmp(264) := "1000" & "000" & "100100110" ;	-- JEQ @Set4
tmp(265) := "1001" & "000" & "000000100" ;	-- CEQ R0, @4
tmp(266) := "1000" & "000" & "100101010" ;	-- JEQ @Set5
tmp(267) := "0101" & "010" & "000000000" ;	-- LDI R2, @0
tmp(268) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(269) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(270) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(271) := "0001" & "101" & "000000000" ;	-- LDA R5, @0
tmp(272) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(273) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(274) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(275) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(276) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(277) := "0110" & "000" & "111111111" ;	-- CLR @KEY0
tmp(278) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(279) := "0110" & "000" & "111111010" ;	-- CLR @SEC
tmp(280) := "1010" & "000" & "001111111" ;	-- JSR @BAS5SET3
tmp(281) := "0111" & "000" & "000101001" ;	-- JMP @Clock

-- LABEL Set1
tmp(282) := "0101" & "010" & "000000010" ;	-- LDI R2, $2
tmp(283) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(284) := "0101" & "000" & "000000001" ;	-- LDI R0, @1
tmp(285) := "0111" & "000" & "010110000" ;	-- JMP @VerificaK0

-- LABEL Set2
tmp(286) := "0101" & "010" & "000000100" ;	-- LDI R2, $4
tmp(287) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(288) := "0101" & "000" & "000000010" ;	-- LDI R0, @2
tmp(289) := "0111" & "000" & "010110000" ;	-- JMP @VerificaK0

-- LABEL Set3
tmp(290) := "0101" & "010" & "000001000" ;	-- LDI R2, $8
tmp(291) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(292) := "0101" & "000" & "000000011" ;	-- LDI R0, @3
tmp(293) := "0111" & "000" & "010110000" ;	-- JMP @VerificaK0

-- LABEL Set4
tmp(294) := "0101" & "010" & "000010000" ;	-- LDI R2, $16
tmp(295) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(296) := "0101" & "000" & "000000100" ;	-- LDI R0, @4
tmp(297) := "0111" & "000" & "010110000" ;	-- JMP @VerificaK0

-- LABEL Set5
tmp(298) := "0101" & "010" & "000100000" ;	-- LDI R2, $32
tmp(299) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(300) := "0101" & "000" & "000000101" ;	-- LDI R0, @5
tmp(301) := "0111" & "000" & "010110000" ;	-- JMP @VerificaK0

		  
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;