library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 16;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant ANDD : std_logic_vector(3 downto 0) := "0100";
  constant LDI  : std_logic_vector(3 downto 0) := "0101";
  constant STA  : std_logic_vector(3 downto 0) := "0110";
  constant JMP  : std_logic_vector(3 downto 0) := "0111";
  constant JEQ  : std_logic_vector(3 downto 0) := "1000";
  constant CEQ  : std_logic_vector(3 downto 0) := "1001";
  constant JSR  : std_logic_vector(3 downto 0) := "1010";
  constant RET  : std_logic_vector(3 downto 0) := "1011";
  constant JNE  : std_logic_vector(3 downto 0) := "1100";
  constant JLT  : std_logic_vector(3 downto 0) := "1101";
  constant CLT  : std_logic_vector(3 downto 0) := "1110";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
  

-- LABEL Setup
tmp(0) := "0101" & "000" & "010000000" ;	-- LDI R0, $128
tmp(1) := "0110" & "000" & "000111111" ;	-- STA @63, R0
tmp(2) := "0101" & "000" & "000000000" ;	-- LDI R0, $0
tmp(3) := "0110" & "000" & "000000000" ;	-- STA @0, R0
tmp(4) := "0101" & "001" & "000000001" ;	-- LDI R1, $1
tmp(5) := "0110" & "001" & "000000001" ;	-- STA @1, R1
tmp(6) := "0101" & "001" & "000000010" ;	-- LDI R1, $2
tmp(7) := "0110" & "001" & "000000010" ;	-- STA @2, R1
tmp(8) := "0101" & "001" & "000000011" ;	-- LDI R1, $3
tmp(9) := "0110" & "001" & "000000011" ;	-- STA @3, R1
tmp(10) := "0110" & "001" & "000011001" ;	-- STA @BAS5, R1
tmp(11) := "0101" & "001" & "000000100" ;	-- LDI R1, $4
tmp(12) := "0110" & "001" & "000000100" ;	-- STA @4, R1
tmp(13) := "0101" & "001" & "000000101" ;	-- LDI R1, $5
tmp(14) := "0110" & "001" & "000000101" ;	-- STA @5, R1
tmp(15) := "0101" & "001" & "000000110" ;	-- LDI R1, $6
tmp(16) := "0110" & "001" & "000000110" ;	-- STA @6, R1
tmp(17) := "0101" & "001" & "000001010" ;	-- LDI R1, $10
tmp(18) := "0110" & "001" & "000001010" ;	-- STA @10, R1
tmp(19) := "0110" & "001" & "000011000" ;	-- STA @BAS4, R1
tmp(20) := "0101" & "001" & "000001001" ;	-- LDI R1, $9
tmp(21) := "0110" & "000" & "000010111" ;	-- STA @FLAG, R0
tmp(22) := "0110" & "001" & "000001011" ;	-- STA @LIM0, R1
tmp(23) := "0110" & "001" & "000001100" ;	-- STA @LIM1, R1
tmp(24) := "0110" & "001" & "000001101" ;	-- STA @LIM2, R1
tmp(25) := "0110" & "001" & "000001110" ;	-- STA @LIM3, R1
tmp(26) := "0110" & "001" & "000001111" ;	-- STA @LIM4, R1
tmp(27) := "0110" & "001" & "000010000" ;	-- STA @LIM5, R1
tmp(28) := "0110" & "000" & "000010001" ;	-- STA @MEM0, R0
tmp(29) := "0110" & "000" & "000010011" ;	-- STA @MEM2, R0
tmp(30) := "0110" & "000" & "000010010" ;	-- STA @MEM1, R0
tmp(31) := "0110" & "000" & "000010100" ;	-- STA @MEM3, R0
tmp(32) := "0110" & "000" & "000010101" ;	-- STA @MEM4, R0
tmp(33) := "0110" & "000" & "000010110" ;	-- STA @MEM5, R0
tmp(34) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(35) := "0110" & "000" & "100100001" ;	-- STA @HEX1, R0
tmp(36) := "0110" & "000" & "100100010" ;	-- STA @HEX2, R0
tmp(37) := "0110" & "000" & "100100011" ;	-- STA @HEX3, R0
tmp(38) := "0110" & "000" & "100100100" ;	-- STA @HEX4, R0
tmp(39) := "0110" & "000" & "100100101" ;	-- STA @HEX5, R0
tmp(40) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(41) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(42) := "0001" & "101" & "000000000" ;	-- LDA R5, @0
tmp(43) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(44) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(45) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(46) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(47) := "0001" & "000" & "000000000" ;	-- LDA R0, @0

-- LABEL Clock
tmp(48) := "0001" & "011" & "000010001" ;	-- LDA R3, @MEM0
tmp(49) := "0110" & "011" & "100100000" ;	-- STA @HEX0, R3
tmp(50) := "0001" & "011" & "000010010" ;	-- LDA R3, @MEM1
tmp(51) := "0110" & "011" & "100100001" ;	-- STA @HEX1, R3
tmp(52) := "0001" & "011" & "000010011" ;	-- LDA R3, @MEM2
tmp(53) := "0110" & "011" & "100100010" ;	-- STA @HEX2, R3
tmp(54) := "0001" & "011" & "000010100" ;	-- LDA R3, @MEM3
tmp(55) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(56) := "0001" & "011" & "000010101" ;	-- LDA R3, @MEM4
tmp(57) := "0110" & "011" & "100100100" ;	-- STA @HEX4, R3
tmp(58) := "0001" & "011" & "000010110" ;	-- LDA R3, @MEM5
tmp(59) := "0110" & "011" & "100100101" ;	-- STA @HEX5, R3
tmp(60) := "0111" & "000" & "000111101" ;	-- JMP @IncClk

-- LABEL IncClk
tmp(61) := "0001" & "111" & "101100101" ;	-- LDA R7, @SEC
tmp(62) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(63) := "1001" & "111" & "000000001" ;	-- CEQ R7, @1
tmp(64) := "1100" & "000" & "010010010" ;	-- JNE @WaitSet
tmp(65) := "0110" & "000" & "111111010" ;	-- CLR @SEC
tmp(66) := "0001" & "000" & "000010001" ;	-- LDA R0, @MEM0
tmp(67) := "0010" & "000" & "000000001" ;	-- SOMA R0, @1
tmp(68) := "1001" & "000" & "000001010" ;	-- CEQ R0, @10
tmp(69) := "1000" & "000" & "001001001" ;	-- JEQ @ResetMem0
tmp(70) := "0110" & "000" & "000010001" ;	-- STA @MEM0, R0
tmp(71) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(72) := "0111" & "000" & "010010010" ;	-- JMP @WaitSet

-- LABEL ResetMem0
tmp(73) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(74) := "0110" & "000" & "000010001" ;	-- STA @MEM0, R0
tmp(75) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(76) := "0001" & "001" & "000010010" ;	-- LDA R1, @MEM1
tmp(77) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(78) := "1001" & "001" & "000000110" ;	-- CEQ R1, @6
tmp(79) := "1000" & "000" & "001010011" ;	-- JEQ @ResetMem1
tmp(80) := "0110" & "001" & "000010010" ;	-- STA @MEM1, R1
tmp(81) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(82) := "0111" & "000" & "010010010" ;	-- JMP @WaitSet

-- LABEL ResetMem1
tmp(83) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(84) := "0110" & "001" & "000010010" ;	-- STA @MEM1, R1
tmp(85) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(86) := "0001" & "010" & "000010011" ;	-- LDA R2, @MEM2
tmp(87) := "0010" & "010" & "000000001" ;	-- SOMA R2, @1
tmp(88) := "1001" & "010" & "000001010" ;	-- CEQ R2, @10
tmp(89) := "1000" & "000" & "001011101" ;	-- JEQ @ResetMem2
tmp(90) := "0110" & "010" & "000010011" ;	-- STA @MEM2, R2
tmp(91) := "0110" & "010" & "100100010" ;	-- STA @HEX2, R2
tmp(92) := "0111" & "000" & "010010010" ;	-- JMP @WaitSet

-- LABEL ResetMem2
tmp(93) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(94) := "0110" & "010" & "000010011" ;	-- STA @MEM2, R2
tmp(95) := "0110" & "010" & "100100010" ;	-- STA @HEX2, R2
tmp(96) := "0001" & "011" & "000010100" ;	-- LDA R3, @MEM3
tmp(97) := "0010" & "011" & "000000001" ;	-- SOMA R3, @1
tmp(98) := "1001" & "011" & "000000110" ;	-- CEQ R3, @6
tmp(99) := "1000" & "000" & "001100111" ;	-- JEQ @ResetMem3
tmp(100) := "0110" & "011" & "000010100" ;	-- STA @MEM3, R3
tmp(101) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(102) := "0111" & "000" & "010010010" ;	-- JMP @WaitSet

-- LABEL ResetMem3
tmp(103) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(104) := "0110" & "011" & "000010100" ;	-- STA @MEM3, R3
tmp(105) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(106) := "0001" & "100" & "000010101" ;	-- LDA R4, @MEM4
tmp(107) := "0010" & "100" & "000000001" ;	-- SOMA R4, @1
tmp(108) := "1001" & "100" & "000011000" ;	-- CEQ R4, @BAS4
tmp(109) := "1000" & "000" & "001110001" ;	-- JEQ @ResetMem4
tmp(110) := "0110" & "100" & "000010101" ;	-- STA @MEM4, R4
tmp(111) := "0110" & "100" & "100100100" ;	-- STA @HEX4, R4
tmp(112) := "0111" & "000" & "010010010" ;	-- JMP @WaitSet

-- LABEL ResetMem4
tmp(113) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(114) := "0110" & "100" & "000010101" ;	-- STA @MEM4, R4
tmp(115) := "0110" & "100" & "100100100" ;	-- STA @HEX4, R4
tmp(116) := "0001" & "101" & "000010110" ;	-- LDA R5, @MEM5
tmp(117) := "0010" & "101" & "000000001" ;	-- SOMA R5, @1
tmp(118) := "1001" & "101" & "000011001" ;	-- CEQ R5, @BAS5
tmp(119) := "1000" & "000" & "010000011" ;	-- JEQ @Zera
tmp(120) := "0110" & "101" & "000010110" ;	-- STA @MEM5, R5
tmp(121) := "0110" & "101" & "100100101" ;	-- STA @HEX5, R5
tmp(122) := "1001" & "101" & "000000010" ;	-- CEQ R5, @2
tmp(123) := "1010" & "000" & "001111101" ;	-- JSR @BAS4SET4
tmp(124) := "0111" & "000" & "010010010" ;	-- JMP @WaitSet

-- LABEL BAS4SET4
tmp(125) := "0101" & "100" & "000000100" ;	-- LDI R4, $4
tmp(126) := "0110" & "100" & "000011000" ;	-- STA @BAS4, R4
tmp(127) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL BAS4SET10
tmp(128) := "0101" & "100" & "000001010" ;	-- LDI R4, $10
tmp(129) := "0110" & "100" & "000011000" ;	-- STA @BAS4, R4
tmp(130) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Zera
tmp(131) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(132) := "0110" & "000" & "000010001" ;	-- STA @MEM0, R0
tmp(133) := "0110" & "000" & "000010011" ;	-- STA @MEM2, R0
tmp(134) := "0110" & "000" & "000010010" ;	-- STA @MEM1, R0
tmp(135) := "0110" & "000" & "000010100" ;	-- STA @MEM3, R0
tmp(136) := "0110" & "000" & "000010101" ;	-- STA @MEM4, R0
tmp(137) := "0110" & "000" & "000010110" ;	-- STA @MEM5, R0
tmp(138) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(139) := "0110" & "000" & "100100001" ;	-- STA @HEX1, R0
tmp(140) := "0110" & "000" & "100100010" ;	-- STA @HEX2, R0
tmp(141) := "0110" & "000" & "100100011" ;	-- STA @HEX3, R0
tmp(142) := "0110" & "000" & "100100100" ;	-- STA @HEX4, R0
tmp(143) := "0110" & "000" & "100100101" ;	-- STA @HEX5, R0
tmp(144) := "1010" & "000" & "010000000" ;	-- JSR @BAS4SET10
tmp(145) := "0111" & "000" & "010010010" ;	-- JMP @WaitSet

-- LABEL WaitSet
tmp(146) := "0001" & "111" & "101100011" ;	-- LDA R7, @KEY3
tmp(147) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(148) := "1001" & "111" & "000000001" ;	-- CEQ R7, @1
tmp(149) := "1000" & "000" & "010010111" ;	-- JEQ @SetMem
tmp(150) := "0111" & "000" & "000111101" ;	-- JMP @IncClk

-- LABEL SetMem
tmp(151) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(152) := "0001" & "011" & "000010001" ;	-- LDA R3, @MEM0
tmp(153) := "0110" & "011" & "100100000" ;	-- STA @HEX0, R3
tmp(154) := "0001" & "011" & "000010010" ;	-- LDA R3, @MEM1
tmp(155) := "0110" & "011" & "100100001" ;	-- STA @HEX1, R3
tmp(156) := "0001" & "011" & "000010011" ;	-- LDA R3, @MEM2
tmp(157) := "0110" & "011" & "100100010" ;	-- STA @HEX2, R3
tmp(158) := "0001" & "011" & "000010100" ;	-- LDA R3, @MEM3
tmp(159) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(160) := "0001" & "011" & "000010101" ;	-- LDA R3, @MEM4
tmp(161) := "0110" & "011" & "100100100" ;	-- STA @HEX4, R3
tmp(162) := "0001" & "011" & "000010110" ;	-- LDA R3, @MEM5
tmp(163) := "0110" & "011" & "100100101" ;	-- STA @HEX5, R3
tmp(164) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(165) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(166) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(167) := "0001" & "010" & "000000001" ;	-- LDA R2, @1
tmp(168) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(169) := "0110" & "000" & "111111111" ;	-- CLR @KEY0
tmp(170) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(171) := "0111" & "000" & "010101100" ;	-- JMP @VerificaK0

-- LABEL VerificaK0
tmp(172) := "0001" & "110" & "101100000" ;	-- LDA R6, @KEY0
tmp(173) := "0100" & "110" & "000000001" ;	-- AND R6, @1
tmp(174) := "1001" & "110" & "000000000" ;	-- CEQ R6, @0
tmp(175) := "1000" & "000" & "010110001" ;	-- JEQ @VerificaK1
tmp(176) := "0111" & "000" & "010110110" ;	-- JMP @IncMem

-- LABEL VerificaK1
tmp(177) := "0001" & "111" & "101100011" ;	-- LDA R7, @KEY3
tmp(178) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(179) := "1001" & "111" & "000000000" ;	-- CEQ R7, @0
tmp(180) := "1100" & "000" & "100000000" ;	-- JNE @Set0
tmp(181) := "0111" & "000" & "010101100" ;	-- JMP @VerificaK0

-- LABEL IncMem
tmp(182) := "0110" & "000" & "111111111" ;	-- CLR @KEY0
tmp(183) := "1001" & "000" & "000000000" ;	-- CEQ R0, @0
tmp(184) := "1000" & "000" & "011000011" ;	-- JEQ @IncMem0
tmp(185) := "1001" & "000" & "000000001" ;	-- CEQ R0, @1
tmp(186) := "1000" & "000" & "011001011" ;	-- JEQ @IncMem1
tmp(187) := "1001" & "000" & "000000010" ;	-- CEQ R0, @2
tmp(188) := "1000" & "000" & "011010011" ;	-- JEQ @IncMem2
tmp(189) := "1001" & "000" & "000000011" ;	-- CEQ R0, @3
tmp(190) := "1000" & "000" & "011011011" ;	-- JEQ @IncMem3
tmp(191) := "1001" & "000" & "000000100" ;	-- CEQ R0, @4
tmp(192) := "1000" & "000" & "011100011" ;	-- JEQ @IncMem4
tmp(193) := "1001" & "000" & "000000101" ;	-- CEQ R0, @5
tmp(194) := "1000" & "000" & "011110010" ;	-- JEQ @IncMem5

-- LABEL IncMem0
tmp(195) := "0001" & "001" & "000010001" ;	-- LDA R1, @MEM0
tmp(196) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(197) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(198) := "1100" & "000" & "011001000" ;	-- JNE @StaMem0
tmp(199) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem0
tmp(200) := "0110" & "001" & "000010001" ;	-- STA @MEM0, R1
tmp(201) := "0110" & "001" & "100100000" ;	-- STA @HEX0, R1
tmp(202) := "0111" & "000" & "010110001" ;	-- JMP @VerificaK1

-- LABEL IncMem1
tmp(203) := "0001" & "001" & "000010010" ;	-- LDA R1, @MEM1
tmp(204) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(205) := "1001" & "001" & "000000110" ;	-- CEQ R1, @6
tmp(206) := "1100" & "000" & "011010000" ;	-- JNE @StaMem1
tmp(207) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem1
tmp(208) := "0110" & "001" & "000010010" ;	-- STA @MEM1, R1
tmp(209) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(210) := "0111" & "000" & "010110001" ;	-- JMP @VerificaK1

-- LABEL IncMem2
tmp(211) := "0001" & "001" & "000010011" ;	-- LDA R1, @MEM2
tmp(212) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(213) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(214) := "1100" & "000" & "011011000" ;	-- JNE @StaMem2
tmp(215) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem2
tmp(216) := "0110" & "001" & "000010011" ;	-- STA @MEM2, R1
tmp(217) := "0110" & "001" & "100100010" ;	-- STA @HEX2, R1
tmp(218) := "0111" & "000" & "010110001" ;	-- JMP @VerificaK1

-- LABEL IncMem3
tmp(219) := "0001" & "001" & "000010100" ;	-- LDA R1, @MEM3
tmp(220) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(221) := "1001" & "001" & "000000110" ;	-- CEQ R1, @6
tmp(222) := "1100" & "000" & "011100000" ;	-- JNE @StaMem3
tmp(223) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem3
tmp(224) := "0110" & "001" & "000010100" ;	-- STA @MEM3, R1
tmp(225) := "0110" & "001" & "100100011" ;	-- STA @HEX3, R1
tmp(226) := "0111" & "000" & "010110001" ;	-- JMP @VerificaK1

-- LABEL IncMem4
tmp(227) := "0001" & "001" & "000010101" ;	-- LDA R1, @MEM4
tmp(228) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(229) := "1001" & "001" & "000011000" ;	-- CEQ R1, @BAS4
tmp(230) := "1100" & "000" & "011101000" ;	-- JNE @StaMem4
tmp(231) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem4
tmp(232) := "0110" & "001" & "000010101" ;	-- STA @MEM4, R1
tmp(233) := "0110" & "001" & "100100100" ;	-- STA @HEX4, R1
tmp(234) := "1110" & "001" & "000000100" ;	-- CLT R1, @4
tmp(235) := "1101" & "000" & "011101111" ;	-- JLT @setMax2
tmp(236) := "0001" & "001" & "000000010" ;	-- LDA R1, @2
tmp(237) := "0110" & "001" & "000011001" ;	-- STA @BAS5, R1
tmp(238) := "0111" & "000" & "010110001" ;	-- JMP @VerificaK1

-- LABEL setMax2
tmp(239) := "0001" & "001" & "000000011" ;	-- LDA R1, @3
tmp(240) := "0110" & "001" & "000011001" ;	-- STA @BAS5, R1
tmp(241) := "0111" & "000" & "010110001" ;	-- JMP @VerificaK1

-- LABEL IncMem5
tmp(242) := "0001" & "001" & "000010110" ;	-- LDA R1, @MEM5
tmp(243) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(244) := "1001" & "001" & "000011001" ;	-- CEQ R1, @BAS5
tmp(245) := "1100" & "000" & "011110111" ;	-- JNE @StaMem5
tmp(246) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaMem5
tmp(247) := "1001" & "001" & "000000010" ;	-- CEQ R1, @2
tmp(248) := "1100" & "000" & "011111011" ;	-- JNE @SetBase24
tmp(249) := "0101" & "001" & "000000100" ;	-- LDI R1, $4
tmp(250) := "0110" & "001" & "000011000" ;	-- STA @BAS4, R1

-- LABEL SetBase24
tmp(251) := "0110" & "001" & "000010110" ;	-- STA @MEM5, R1
tmp(252) := "0110" & "001" & "100100101" ;	-- STA @HEX5, R1
tmp(253) := "0001" & "001" & "000000011" ;	-- LDA R1, @3
tmp(254) := "0110" & "001" & "000011001" ;	-- STA @BAS5, R1
tmp(255) := "0111" & "000" & "010110001" ;	-- JMP @VerificaK1

-- LABEL Set0
tmp(256) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(257) := "1001" & "000" & "000000000" ;	-- CEQ R0, @0
tmp(258) := "1000" & "000" & "100011001" ;	-- JEQ @Set1
tmp(259) := "1001" & "000" & "000000001" ;	-- CEQ R0, @1
tmp(260) := "1000" & "000" & "100011101" ;	-- JEQ @Set2
tmp(261) := "1001" & "000" & "000000010" ;	-- CEQ R0, @2
tmp(262) := "1000" & "000" & "100100001" ;	-- JEQ @Set3
tmp(263) := "1001" & "000" & "000000011" ;	-- CEQ R0, @3
tmp(264) := "1000" & "000" & "100100101" ;	-- JEQ @Set4
tmp(265) := "1001" & "000" & "000000100" ;	-- CEQ R0, @4
tmp(266) := "1000" & "000" & "100101001" ;	-- JEQ @Set5
tmp(267) := "0101" & "010" & "000000000" ;	-- LDI R2, @0
tmp(268) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(269) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(270) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(271) := "0001" & "101" & "000000000" ;	-- LDA R5, @0
tmp(272) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(273) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(274) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(275) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(276) := "0001" & "000" & "000000000" ;	-- LDA R0, @0
tmp(277) := "0110" & "000" & "111111111" ;	-- CLR @KEY0
tmp(278) := "0110" & "000" & "111111100" ;	-- CLR @KEY3
tmp(279) := "0110" & "000" & "000010111" ;	-- STA @FLAG, R0
tmp(280) := "0111" & "000" & "000110000" ;	-- JMP @Clock

-- LABEL Set1
tmp(281) := "0101" & "010" & "000000010" ;	-- LDI R2, $2
tmp(282) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(283) := "0101" & "000" & "000000001" ;	-- LDI R0, @1
tmp(284) := "0111" & "000" & "010101100" ;	-- JMP @VerificaK0

-- LABEL Set2
tmp(285) := "0101" & "010" & "000000100" ;	-- LDI R2, $4
tmp(286) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(287) := "0101" & "000" & "000000010" ;	-- LDI R0, @2
tmp(288) := "0111" & "000" & "010101100" ;	-- JMP @VerificaK0

-- LABEL Set3
tmp(289) := "0101" & "010" & "000001000" ;	-- LDI R2, $8
tmp(290) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(291) := "0101" & "000" & "000000011" ;	-- LDI R0, @3
tmp(292) := "0111" & "000" & "010101100" ;	-- JMP @VerificaK0

-- LABEL Set4
tmp(293) := "0101" & "010" & "000010000" ;	-- LDI R2, $16
tmp(294) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(295) := "0101" & "000" & "000000100" ;	-- LDI R0, @4
tmp(296) := "0111" & "000" & "010101100" ;	-- JMP @VerificaK0

-- LABEL Set5
tmp(297) := "0101" & "010" & "000100000" ;	-- LDI R2, $32
tmp(298) := "0110" & "010" & "100000000" ;	-- STA @LEDb, R2
tmp(299) := "0101" & "000" & "000000101" ;	-- LDI R0, @5
tmp(300) := "0111" & "000" & "010101100" ;	-- JMP @VerificaK0

		  
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;