library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 16;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant ANDD : std_logic_vector(3 downto 0) := "0100";
  constant LDI  : std_logic_vector(3 downto 0) := "0101";
  constant STA  : std_logic_vector(3 downto 0) := "0110";
  constant JMP  : std_logic_vector(3 downto 0) := "0111";
  constant JEQ  : std_logic_vector(3 downto 0) := "1000";
  constant CEQ  : std_logic_vector(3 downto 0) := "1001";
  constant JSR  : std_logic_vector(3 downto 0) := "1010";
  constant RET  : std_logic_vector(3 downto 0) := "1011";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
  

-- LABEL Setup
tmp(0) := "0101" & "000" & "000000000" ;	-- LDI R0, $0
tmp(1) := "0110" & "000" & "000000000" ;	-- STA @0, R0
tmp(2) := "0101" & "001" & "000000001" ;	-- LDI R1, $1
tmp(3) := "0110" & "001" & "000000001" ;	-- STA @1, R1
tmp(4) := "0101" & "001" & "000000010" ;	-- LDI R1, $2
tmp(5) := "0110" & "001" & "000000010" ;	-- STA @2, R1
tmp(6) := "0101" & "001" & "000000011" ;	-- LDI R1, $3
tmp(7) := "0110" & "001" & "000000011" ;	-- STA @3, R1
tmp(8) := "0101" & "001" & "000000100" ;	-- LDI R1, $4
tmp(9) := "0110" & "001" & "000000100" ;	-- STA @4, R1
tmp(10) := "0101" & "001" & "000000101" ;	-- LDI R1, $5
tmp(11) := "0110" & "001" & "000000101" ;	-- STA @5, R1
tmp(12) := "0101" & "001" & "000001010" ;	-- LDI R1, $10
tmp(13) := "0110" & "001" & "000001010" ;	-- STA @10, R1
tmp(14) := "0110" & "000" & "000010011" ;	-- STA @FLAG, R0
tmp(15) := "0110" & "000" & "000000110" ;	-- STA @LIM0, R0
tmp(16) := "0110" & "000" & "000000111" ;	-- STA @LIM1, R0
tmp(17) := "0110" & "000" & "000001000" ;	-- STA @LIM2, R0
tmp(18) := "0110" & "000" & "000001001" ;	-- STA @LIM3, R0
tmp(19) := "0110" & "000" & "000001011" ;	-- STA @LIM4, R0
tmp(20) := "0110" & "000" & "000001100" ;	-- STA @LIM5, R0
tmp(21) := "0110" & "000" & "000001101" ;	-- STA @MEM0, R0
tmp(22) := "0110" & "000" & "000001110" ;	-- STA @MEM1, R0
tmp(23) := "0110" & "000" & "000001111" ;	-- STA @MEM2, R0
tmp(24) := "0110" & "000" & "000010000" ;	-- STA @MEM3, R0
tmp(25) := "0110" & "000" & "000010001" ;	-- STA @MEM4, R0
tmp(26) := "0110" & "000" & "000010010" ;	-- STA @MEM5, R0
tmp(27) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(28) := "0110" & "000" & "100100001" ;	-- STA @HEX1, R0
tmp(29) := "0110" & "000" & "100100010" ;	-- STA @HEX2, R0
tmp(30) := "0110" & "000" & "100100011" ;	-- STA @HEX3, R0
tmp(31) := "0110" & "000" & "100100100" ;	-- STA @HEX4, R0
tmp(32) := "0110" & "000" & "100100101" ;	-- STA @HEX5, R0
tmp(33) := "0001" & "111" & "000000000" ;	-- LDA R7, @0
tmp(34) := "0001" & "110" & "000000000" ;	-- LDA R6, @0
tmp(35) := "0001" & "101" & "000000000" ;	-- LDA R5, @0
tmp(36) := "0001" & "100" & "000000000" ;	-- LDA R4, @0
tmp(37) := "0001" & "011" & "000000000" ;	-- LDA R3, @0
tmp(38) := "0001" & "010" & "000000000" ;	-- LDA R2, @0
tmp(39) := "0001" & "001" & "000000000" ;	-- LDA R1, @0
tmp(40) := "0001" & "000" & "000000000" ;	-- LDA R0, @0

-- LABEL VerificaK0
tmp(41) := "0001" & "110" & "101100000" ;	-- LDA R6, @KEY0
tmp(42) := "0100" & "110" & "000000001" ;	-- AND R6, @1
tmp(43) := "1001" & "110" & "000000000" ;	-- CEQ R6, @0
tmp(44) := "1000" & "000" & "000101110" ;	-- JEQ @VerificaK1
tmp(45) := "1010" & "000" & "000110100" ;	-- JSR @IncLim

-- LABEL VerificaK1
tmp(46) := "0001" & "111" & "101100001" ;	-- LDA R7, @KEY1
tmp(47) := "0100" & "111" & "000000001" ;	-- AND R7, @1
tmp(48) := "1001" & "111" & "000000000" ;	-- CEQ R7, @0
tmp(49) := "1000" & "000" & "000101001" ;	-- JEQ @VerificaK0
tmp(50) := "1010" & "000" & "001110111" ;	-- JSR @Set0
tmp(51) := "0111" & "000" & "000101001" ;	-- JMP @VerificaK0

-- LABEL IncLim
tmp(52) := "0110" & "000" & "111111111" ;	-- CLR @KEY0
tmp(53) := "1001" & "000" & "000000000" ;	-- CEQ R0, @0
tmp(54) := "1000" & "000" & "001000001" ;	-- JEQ @IncLim0
tmp(55) := "1001" & "000" & "000000001" ;	-- CEQ R0, @1
tmp(56) := "1000" & "000" & "001001010" ;	-- JEQ @IncLim1
tmp(57) := "1001" & "000" & "000000010" ;	-- CEQ R0, @2
tmp(58) := "1000" & "000" & "001010011" ;	-- JEQ @IncLim2
tmp(59) := "1001" & "000" & "000000011" ;	-- CEQ R0, @3
tmp(60) := "1000" & "000" & "001011100" ;	-- JEQ @IncLim3
tmp(61) := "1001" & "000" & "000000100" ;	-- CEQ R0, @4
tmp(62) := "1000" & "000" & "001100101" ;	-- JEQ @IncLim4
tmp(63) := "1001" & "000" & "000000101" ;	-- CEQ R0, @5
tmp(64) := "1000" & "000" & "001101110" ;	-- JEQ @IncLim5

-- LABEL IncLim0
tmp(65) := "0001" & "001" & "000000110" ;	-- LDA R1, @LIM0
tmp(66) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(67) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(68) := "1000" & "000" & "001000110" ;	-- JEQ @ResetLim0
tmp(69) := "0111" & "000" & "001000111" ;	-- JMP @StaLim0

-- LABEL ResetLim0
tmp(70) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaLim0
tmp(71) := "0110" & "001" & "000000110" ;	-- STA @LIM0, R1
tmp(72) := "0110" & "001" & "100100000" ;	-- STA @HEX0, R1
tmp(73) := "0111" & "000" & "000101110" ;	-- JMP @VerificaK1

-- LABEL IncLim1
tmp(74) := "0001" & "001" & "000000111" ;	-- LDA R1, @LIM1
tmp(75) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(76) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(77) := "1000" & "000" & "001001111" ;	-- JEQ @ResetLim1
tmp(78) := "0111" & "000" & "001010000" ;	-- JMP @StaLim1

-- LABEL ResetLim1
tmp(79) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaLim1
tmp(80) := "0110" & "001" & "000000111" ;	-- STA @LIM1, R1
tmp(81) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(82) := "0111" & "000" & "000101110" ;	-- JMP @VerificaK1

-- LABEL IncLim2
tmp(83) := "0001" & "001" & "000001000" ;	-- LDA R1, @LIM2
tmp(84) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(85) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(86) := "1000" & "000" & "001011000" ;	-- JEQ @ResetLim2
tmp(87) := "0111" & "000" & "001011001" ;	-- JMP @StaLim2

-- LABEL ResetLim2
tmp(88) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaLim2
tmp(89) := "0110" & "001" & "000001000" ;	-- STA @LIM2, R1
tmp(90) := "0110" & "001" & "100100010" ;	-- STA @HEX2, R1
tmp(91) := "0111" & "000" & "000101110" ;	-- JMP @VerificaK1

-- LABEL IncLim3
tmp(92) := "0001" & "001" & "000001001" ;	-- LDA R1, @LIM3
tmp(93) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(94) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(95) := "1000" & "000" & "001100001" ;	-- JEQ @ResetLim3
tmp(96) := "0111" & "000" & "001100010" ;	-- JMP @StaLim3

-- LABEL ResetLim3
tmp(97) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaLim3
tmp(98) := "0110" & "001" & "000001001" ;	-- STA @LIM3, R1
tmp(99) := "0110" & "001" & "100100011" ;	-- STA @HEX3, R1
tmp(100) := "0111" & "000" & "000101110" ;	-- JMP @VerificaK1

-- LABEL IncLim4
tmp(101) := "0001" & "001" & "000001011" ;	-- LDA R1, @LIM4
tmp(102) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(103) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(104) := "1000" & "000" & "001101010" ;	-- JEQ @ResetLim4
tmp(105) := "0111" & "000" & "001101011" ;	-- JMP @StaLim4

-- LABEL ResetLim4
tmp(106) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaLim4
tmp(107) := "0110" & "001" & "000001011" ;	-- STA @LIM4, R1
tmp(108) := "0110" & "001" & "100100100" ;	-- STA @HEX4, R1
tmp(109) := "0111" & "000" & "000101110" ;	-- JMP @VerificaK1

-- LABEL IncLim5
tmp(110) := "0001" & "001" & "000001100" ;	-- LDA R1, @LIM5
tmp(111) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(112) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(113) := "1000" & "000" & "001110011" ;	-- JEQ @ResetLim5
tmp(114) := "0111" & "000" & "001110100" ;	-- JMP @StaLim5

-- LABEL ResetLim5
tmp(115) := "0001" & "001" & "000000000" ;	-- LDA R1, $0

-- LABEL StaLim5
tmp(116) := "0110" & "001" & "000001100" ;	-- STA @LIM5, R1
tmp(117) := "0110" & "001" & "100100101" ;	-- STA @HEX5, R1
tmp(118) := "0111" & "000" & "000101110" ;	-- JMP @VerificaK1

-- LABEL Set0
tmp(119) := "0110" & "000" & "111111110" ;	-- CLR @KEY1
tmp(120) := "1001" & "000" & "000000000" ;	-- CEQ R0, @0
tmp(121) := "1000" & "000" & "010000011" ;	-- JEQ @Set1
tmp(122) := "1001" & "000" & "000000001" ;	-- CEQ R0, @1
tmp(123) := "1000" & "000" & "010000101" ;	-- JEQ @Set2
tmp(124) := "1001" & "000" & "000000010" ;	-- CEQ R0, @2
tmp(125) := "1000" & "000" & "010000111" ;	-- JEQ @Set3
tmp(126) := "1001" & "000" & "000000011" ;	-- CEQ R0, @3
tmp(127) := "1000" & "000" & "010001001" ;	-- JEQ @Set4
tmp(128) := "1001" & "000" & "000000100" ;	-- CEQ R0, @4
tmp(129) := "1000" & "000" & "010001011" ;	-- JEQ @Set5
tmp(130) := "0111" & "000" & "010001101" ;	-- JMP @Contador

-- LABEL Set1
tmp(131) := "0101" & "000" & "000000001" ;	-- LDI R0, @1
tmp(132) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Set2
tmp(133) := "0101" & "000" & "000000010" ;	-- LDI R0, @2
tmp(134) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Set3
tmp(135) := "0101" & "000" & "000000011" ;	-- LDI R0, @3
tmp(136) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Set4
tmp(137) := "0101" & "000" & "000000100" ;	-- LDI R0, @4
tmp(138) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Set5
tmp(139) := "0101" & "000" & "000000101" ;	-- LDI R0, @5
tmp(140) := "1011" & "000" & "000000000" ;	-- RET

-- LABEL Contador
tmp(141) := "0001" & "011" & "000000001" ;	-- LDA R3, @1
tmp(142) := "0110" & "011" & "100000010" ;	-- STA @LED9, R3
tmp(143) := "0110" & "011" & "100100000" ;	-- STA @HEX0, R3
tmp(144) := "0110" & "011" & "100100001" ;	-- STA @HEX1, R3
tmp(145) := "0110" & "011" & "100100010" ;	-- STA @HEX2, R3
tmp(146) := "0110" & "011" & "100100011" ;	-- STA @HEX3, R3
tmp(147) := "0110" & "011" & "100100100" ;	-- STA @HEX4, R3
tmp(148) := "0110" & "011" & "100100101" ;	-- STA @HEX5, R3
tmp(149) := "0111" & "000" & "010001101" ;	-- JMP @Contador

-- LABEL VerificaK2
tmp(150) := "0001" & "110" & "101100010" ;	-- LDA R6, @KEY2
tmp(151) := "0100" & "110" & "000000001" ;	-- AND R6, @1
tmp(152) := "1001" & "110" & "000000001" ;	-- CEQ R6, @1
tmp(153) := "1000" & "000" & "010011011" ;	-- JEQ @IncMem0
tmp(154) := "0111" & "000" & "010010110" ;	-- JMP @VerificaK2

-- LABEL IncMem0
tmp(155) := "0001" & "000" & "000001101" ;	-- LDA R0, @MEM0
tmp(156) := "0010" & "000" & "000000001" ;	-- SOMA R0, @1
tmp(157) := "1001" & "000" & "000001010" ;	-- CEQ R0, @10
tmp(158) := "1000" & "000" & "010100010" ;	-- JEQ @ResetMem0
tmp(159) := "0110" & "000" & "000001101" ;	-- STA @MEM0, R0
tmp(160) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(161) := "0111" & "000" & "010010110" ;	-- JMP @VerificaK2

-- LABEL ResetMem0
tmp(162) := "0001" & "000" & "000000000" ;	-- LDA R0, $0
tmp(163) := "0110" & "000" & "100100000" ;	-- STA @HEX0, R0
tmp(164) := "0001" & "001" & "000001110" ;	-- LDA R1, @MEM1
tmp(165) := "0010" & "001" & "000000001" ;	-- SOMA R1, @1
tmp(166) := "1001" & "001" & "000001010" ;	-- CEQ R1, @10
tmp(167) := "1000" & "000" & "000000000" ;	-- JEQ ResetMem1
tmp(168) := "0110" & "001" & "000001110" ;	-- STA @MEM1, R1
tmp(169) := "0110" & "001" & "100100001" ;	-- STA @HEX1, R1
tmp(170) := "0111" & "000" & "010010110" ;	-- JMP @VerificaK2

-- LABEL ResetMem1
tmp(171) := "0111" & "000" & "010010110" ;	-- JMP @VerificaK2

		  
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;